-- ======================================================
-- ROM generada autom�ticamente con Python
-- Fecha: 2026-01-13 20:33:31
-- Tama�o: 16384 bytes
-- Ancho de datos: 8 bits
-- Ancho de direcci�n: 14 bits
-- Offset inicial: 0
-- ======================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY rom IS
    port (
    clk      : in  std_logic;
    address  : in  std_logic_vector(13 downto 0);
    data_out : out std_logic_vector(7 downto 0)
    );
END entity;

architecture rtl of rom is
BEGIN

	PROCESS(clk)

    variable addr : std_logic_vector(15 downto 0);

	BEGIN
    if rising_edge(clk) then
        addr:="00"&address;
        case addr is

            when x"0000" => data_out<= x"A2";
        when x"0001" => data_out<= x"FF";
        when x"0002" => data_out<= x"9A";
        when x"0003" => data_out<= x"A9";
        when x"0004" => data_out<= x"FF";
        when x"0005" => data_out<= x"85";
        when x"0006" => data_out<= x"0C";
        when x"0007" => data_out<= x"A9";
        when x"0008" => data_out<= x"3F";
        when x"0009" => data_out<= x"85";
        when x"000A" => data_out<= x"0D";
        when x"000B" => data_out<= x"20";
        when x"000C" => data_out<= x"17";
        when x"000D" => data_out<= x"80";
        when x"000E" => data_out<= x"20";
        when x"000F" => data_out<= x"63";
        when x"0010" => data_out<= x"80";
        when x"0011" => data_out<= x"20";
        when x"0012" => data_out<= x"A4";
        when x"0013" => data_out<= x"80";
        when x"0014" => data_out<= x"4C";
        when x"0015" => data_out<= x"14";
        when x"0016" => data_out<= x"80";
        when x"0017" => data_out<= x"A9";
        when x"0018" => data_out<= x"06";
        when x"0019" => data_out<= x"09";
        when x"001A" => data_out<= x"00";
        when x"001B" => data_out<= x"F0";
        when x"001C" => data_out<= x"45";
        when x"001D" => data_out<= x"A9";
        when x"001E" => data_out<= x"85";
        when x"001F" => data_out<= x"8D";
        when x"0020" => data_out<= x"02";
        when x"0021" => data_out<= x"00";
        when x"0022" => data_out<= x"A9";
        when x"0023" => data_out<= x"BD";
        when x"0024" => data_out<= x"8D";
        when x"0025" => data_out<= x"03";
        when x"0026" => data_out<= x"00";
        when x"0027" => data_out<= x"A9";
        when x"0028" => data_out<= x"00";
        when x"0029" => data_out<= x"8D";
        when x"002A" => data_out<= x"04";
        when x"002B" => data_out<= x"00";
        when x"002C" => data_out<= x"A9";
        when x"002D" => data_out<= x"02";
        when x"002E" => data_out<= x"8D";
        when x"002F" => data_out<= x"05";
        when x"0030" => data_out<= x"00";
        when x"0031" => data_out<= x"A9";
        when x"0032" => data_out<= x"06";
        when x"0033" => data_out<= x"8D";
        when x"0034" => data_out<= x"06";
        when x"0035" => data_out<= x"00";
        when x"0036" => data_out<= x"A9";
        when x"0037" => data_out<= x"00";
        when x"0038" => data_out<= x"8D";
        when x"0039" => data_out<= x"07";
        when x"003A" => data_out<= x"00";
        when x"003B" => data_out<= x"A0";
        when x"003C" => data_out<= x"00";
        when x"003D" => data_out<= x"B1";
        when x"003E" => data_out<= x"02";
        when x"003F" => data_out<= x"91";
        when x"0040" => data_out<= x"04";
        when x"0041" => data_out<= x"C8";
        when x"0042" => data_out<= x"D0";
        when x"0043" => data_out<= x"06";
        when x"0044" => data_out<= x"EE";
        when x"0045" => data_out<= x"03";
        when x"0046" => data_out<= x"00";
        when x"0047" => data_out<= x"EE";
        when x"0048" => data_out<= x"05";
        when x"0049" => data_out<= x"00";
        when x"004A" => data_out<= x"AD";
        when x"004B" => data_out<= x"06";
        when x"004C" => data_out<= x"00";
        when x"004D" => data_out<= x"D0";
        when x"004E" => data_out<= x"08";
        when x"004F" => data_out<= x"AD";
        when x"0050" => data_out<= x"07";
        when x"0051" => data_out<= x"00";
        when x"0052" => data_out<= x"F0";
        when x"0053" => data_out<= x"0E";
        when x"0054" => data_out<= x"CE";
        when x"0055" => data_out<= x"07";
        when x"0056" => data_out<= x"00";
        when x"0057" => data_out<= x"CE";
        when x"0058" => data_out<= x"06";
        when x"0059" => data_out<= x"00";
        when x"005A" => data_out<= x"AD";
        when x"005B" => data_out<= x"06";
        when x"005C" => data_out<= x"00";
        when x"005D" => data_out<= x"0D";
        when x"005E" => data_out<= x"07";
        when x"005F" => data_out<= x"00";
        when x"0060" => data_out<= x"D0";
        when x"0061" => data_out<= x"DB";
        when x"0062" => data_out<= x"60";
        when x"0063" => data_out<= x"A9";
        when x"0064" => data_out<= x"4E";
        when x"0065" => data_out<= x"09";
        when x"0066" => data_out<= x"04";
        when x"0067" => data_out<= x"F0";
        when x"0068" => data_out<= x"3A";
        when x"0069" => data_out<= x"A9";
        when x"006A" => data_out<= x"06";
        when x"006B" => data_out<= x"8D";
        when x"006C" => data_out<= x"02";
        when x"006D" => data_out<= x"00";
        when x"006E" => data_out<= x"A9";
        when x"006F" => data_out<= x"02";
        when x"0070" => data_out<= x"8D";
        when x"0071" => data_out<= x"03";
        when x"0072" => data_out<= x"00";
        when x"0073" => data_out<= x"A9";
        when x"0074" => data_out<= x"4E";
        when x"0075" => data_out<= x"8D";
        when x"0076" => data_out<= x"06";
        when x"0077" => data_out<= x"00";
        when x"0078" => data_out<= x"A9";
        when x"0079" => data_out<= x"04";
        when x"007A" => data_out<= x"8D";
        when x"007B" => data_out<= x"07";
        when x"007C" => data_out<= x"00";
        when x"007D" => data_out<= x"A0";
        when x"007E" => data_out<= x"00";
        when x"007F" => data_out<= x"A9";
        when x"0080" => data_out<= x"00";
        when x"0081" => data_out<= x"91";
        when x"0082" => data_out<= x"02";
        when x"0083" => data_out<= x"C8";
        when x"0084" => data_out<= x"D0";
        when x"0085" => data_out<= x"03";
        when x"0086" => data_out<= x"EE";
        when x"0087" => data_out<= x"03";
        when x"0088" => data_out<= x"00";
        when x"0089" => data_out<= x"AE";
        when x"008A" => data_out<= x"06";
        when x"008B" => data_out<= x"00";
        when x"008C" => data_out<= x"D0";
        when x"008D" => data_out<= x"08";
        when x"008E" => data_out<= x"AE";
        when x"008F" => data_out<= x"07";
        when x"0090" => data_out<= x"00";
        when x"0091" => data_out<= x"F0";
        when x"0092" => data_out<= x"10";
        when x"0093" => data_out<= x"CE";
        when x"0094" => data_out<= x"07";
        when x"0095" => data_out<= x"00";
        when x"0096" => data_out<= x"CE";
        when x"0097" => data_out<= x"06";
        when x"0098" => data_out<= x"00";
        when x"0099" => data_out<= x"AE";
        when x"009A" => data_out<= x"06";
        when x"009B" => data_out<= x"00";
        when x"009C" => data_out<= x"D0";
        when x"009D" => data_out<= x"E3";
        when x"009E" => data_out<= x"AE";
        when x"009F" => data_out<= x"07";
        when x"00A0" => data_out<= x"00";
        when x"00A1" => data_out<= x"D0";
        when x"00A2" => data_out<= x"DE";
        when x"00A3" => data_out<= x"60";
        when x"00A4" => data_out<= x"A2";
        when x"00A5" => data_out<= x"00";
        when x"00A6" => data_out<= x"A9";
        when x"00A7" => data_out<= x"C0";
        when x"00A8" => data_out<= x"8D";
        when x"00A9" => data_out<= x"03";
        when x"00AA" => data_out<= x"C0";
        when x"00AB" => data_out<= x"A2";
        when x"00AC" => data_out<= x"00";
        when x"00AD" => data_out<= x"A9";
        when x"00AE" => data_out<= x"00";
        when x"00AF" => data_out<= x"8D";
        when x"00B0" => data_out<= x"01";
        when x"00B1" => data_out<= x"C0";
        when x"00B2" => data_out<= x"20";
        when x"00B3" => data_out<= x"E5";
        when x"00B4" => data_out<= x"80";
        when x"00B5" => data_out<= x"A9";
        when x"00B6" => data_out<= x"9D";
        when x"00B7" => data_out<= x"A2";
        when x"00B8" => data_out<= x"B1";
        when x"00B9" => data_out<= x"20";
        when x"00BA" => data_out<= x"22";
        when x"00BB" => data_out<= x"81";
        when x"00BC" => data_out<= x"A9";
        when x"00BD" => data_out<= x"80";
        when x"00BE" => data_out<= x"A2";
        when x"00BF" => data_out<= x"B1";
        when x"00C0" => data_out<= x"20";
        when x"00C1" => data_out<= x"22";
        when x"00C2" => data_out<= x"81";
        when x"00C3" => data_out<= x"A9";
        when x"00C4" => data_out<= x"B9";
        when x"00C5" => data_out<= x"A2";
        when x"00C6" => data_out<= x"B1";
        when x"00C7" => data_out<= x"20";
        when x"00C8" => data_out<= x"22";
        when x"00C9" => data_out<= x"81";
        when x"00CA" => data_out<= x"20";
        when x"00CB" => data_out<= x"4E";
        when x"00CC" => data_out<= x"81";
        when x"00CD" => data_out<= x"4C";
        when x"00CE" => data_out<= x"DA";
        when x"00CF" => data_out<= x"80";
        when x"00D0" => data_out<= x"20";
        when x"00D1" => data_out<= x"5C";
        when x"00D2" => data_out<= x"81";
        when x"00D3" => data_out<= x"A9";
        when x"00D4" => data_out<= x"A0";
        when x"00D5" => data_out<= x"A2";
        when x"00D6" => data_out<= x"B1";
        when x"00D7" => data_out<= x"20";
        when x"00D8" => data_out<= x"22";
        when x"00D9" => data_out<= x"81";
        when x"00DA" => data_out<= x"4C";
        when x"00DB" => data_out<= x"D0";
        when x"00DC" => data_out<= x"80";
        when x"00DD" => data_out<= x"A2";
        when x"00DE" => data_out<= x"00";
        when x"00DF" => data_out<= x"A9";
        when x"00E0" => data_out<= x"00";
        when x"00E1" => data_out<= x"4C";
        when x"00E2" => data_out<= x"E4";
        when x"00E3" => data_out<= x"80";
        when x"00E4" => data_out<= x"60";
        when x"00E5" => data_out<= x"A9";
        when x"00E6" => data_out<= x"80";
        when x"00E7" => data_out<= x"8D";
        when x"00E8" => data_out<= x"21";
        when x"00E9" => data_out<= x"C0";
        when x"00EA" => data_out<= x"A9";
        when x"00EB" => data_out<= x"00";
        when x"00EC" => data_out<= x"8D";
        when x"00ED" => data_out<= x"21";
        when x"00EE" => data_out<= x"C0";
        when x"00EF" => data_out<= x"60";
        when x"00F0" => data_out<= x"48";
        when x"00F1" => data_out<= x"AD";
        when x"00F2" => data_out<= x"21";
        when x"00F3" => data_out<= x"C0";
        when x"00F4" => data_out<= x"29";
        when x"00F5" => data_out<= x"01";
        when x"00F6" => data_out<= x"F0";
        when x"00F7" => data_out<= x"F9";
        when x"00F8" => data_out<= x"68";
        when x"00F9" => data_out<= x"8D";
        when x"00FA" => data_out<= x"20";
        when x"00FB" => data_out<= x"C0";
        when x"00FC" => data_out<= x"60";
        when x"00FD" => data_out<= x"AD";
        when x"00FE" => data_out<= x"21";
        when x"00FF" => data_out<= x"C0";
        when x"0100" => data_out<= x"29";
        when x"0101" => data_out<= x"02";
        when x"0102" => data_out<= x"F0";
        when x"0103" => data_out<= x"F9";
        when x"0104" => data_out<= x"AD";
        when x"0105" => data_out<= x"20";
        when x"0106" => data_out<= x"C0";
        when x"0107" => data_out<= x"A2";
        when x"0108" => data_out<= x"00";
        when x"0109" => data_out<= x"60";
        when x"010A" => data_out<= x"AD";
        when x"010B" => data_out<= x"21";
        when x"010C" => data_out<= x"C0";
        when x"010D" => data_out<= x"29";
        when x"010E" => data_out<= x"02";
        when x"010F" => data_out<= x"F0";
        when x"0110" => data_out<= x"02";
        when x"0111" => data_out<= x"A9";
        when x"0112" => data_out<= x"01";
        when x"0113" => data_out<= x"A2";
        when x"0114" => data_out<= x"00";
        when x"0115" => data_out<= x"60";
        when x"0116" => data_out<= x"AD";
        when x"0117" => data_out<= x"21";
        when x"0118" => data_out<= x"C0";
        when x"0119" => data_out<= x"29";
        when x"011A" => data_out<= x"01";
        when x"011B" => data_out<= x"F0";
        when x"011C" => data_out<= x"02";
        when x"011D" => data_out<= x"A9";
        when x"011E" => data_out<= x"01";
        when x"011F" => data_out<= x"A2";
        when x"0120" => data_out<= x"00";
        when x"0121" => data_out<= x"60";
        when x"0122" => data_out<= x"8D";
        when x"0123" => data_out<= x"14";
        when x"0124" => data_out<= x"00";
        when x"0125" => data_out<= x"8E";
        when x"0126" => data_out<= x"15";
        when x"0127" => data_out<= x"00";
        when x"0128" => data_out<= x"A0";
        when x"0129" => data_out<= x"00";
        when x"012A" => data_out<= x"B1";
        when x"012B" => data_out<= x"14";
        when x"012C" => data_out<= x"F0";
        when x"012D" => data_out<= x"14";
        when x"012E" => data_out<= x"48";
        when x"012F" => data_out<= x"AD";
        when x"0130" => data_out<= x"21";
        when x"0131" => data_out<= x"C0";
        when x"0132" => data_out<= x"29";
        when x"0133" => data_out<= x"01";
        when x"0134" => data_out<= x"F0";
        when x"0135" => data_out<= x"F9";
        when x"0136" => data_out<= x"68";
        when x"0137" => data_out<= x"8D";
        when x"0138" => data_out<= x"20";
        when x"0139" => data_out<= x"C0";
        when x"013A" => data_out<= x"C8";
        when x"013B" => data_out<= x"D0";
        when x"013C" => data_out<= x"ED";
        when x"013D" => data_out<= x"EE";
        when x"013E" => data_out<= x"15";
        when x"013F" => data_out<= x"00";
        when x"0140" => data_out<= x"D0";
        when x"0141" => data_out<= x"E8";
        when x"0142" => data_out<= x"60";
        when x"0143" => data_out<= x"A9";
        when x"0144" => data_out<= x"80";
        when x"0145" => data_out<= x"8D";
        when x"0146" => data_out<= x"21";
        when x"0147" => data_out<= x"C0";
        when x"0148" => data_out<= x"A9";
        when x"0149" => data_out<= x"00";
        when x"014A" => data_out<= x"8D";
        when x"014B" => data_out<= x"21";
        when x"014C" => data_out<= x"C0";
        when x"014D" => data_out<= x"60";
        when x"014E" => data_out<= x"A9";
        when x"014F" => data_out<= x"00";
        when x"0150" => data_out<= x"8D";
        when x"0151" => data_out<= x"46";
        when x"0152" => data_out<= x"02";
        when x"0153" => data_out<= x"A2";
        when x"0154" => data_out<= x"02";
        when x"0155" => data_out<= x"8D";
        when x"0156" => data_out<= x"00";
        when x"0157" => data_out<= x"02";
        when x"0158" => data_out<= x"8E";
        when x"0159" => data_out<= x"01";
        when x"015A" => data_out<= x"02";
        when x"015B" => data_out<= x"60";
        when x"015C" => data_out<= x"20";
        when x"015D" => data_out<= x"6A";
        when x"015E" => data_out<= x"AE";
        when x"015F" => data_out<= x"A9";
        when x"0160" => data_out<= x"FF";
        when x"0161" => data_out<= x"8D";
        when x"0162" => data_out<= x"01";
        when x"0163" => data_out<= x"C0";
        when x"0164" => data_out<= x"20";
        when x"0165" => data_out<= x"45";
        when x"0166" => data_out<= x"8C";
        when x"0167" => data_out<= x"A9";
        when x"0168" => data_out<= x"93";
        when x"0169" => data_out<= x"A2";
        when x"016A" => data_out<= x"B3";
        when x"016B" => data_out<= x"20";
        when x"016C" => data_out<= x"22";
        when x"016D" => data_out<= x"81";
        when x"016E" => data_out<= x"20";
        when x"016F" => data_out<= x"45";
        when x"0170" => data_out<= x"8C";
        when x"0171" => data_out<= x"A9";
        when x"0172" => data_out<= x"27";
        when x"0173" => data_out<= x"A2";
        when x"0174" => data_out<= x"B6";
        when x"0175" => data_out<= x"20";
        when x"0176" => data_out<= x"22";
        when x"0177" => data_out<= x"81";
        when x"0178" => data_out<= x"20";
        when x"0179" => data_out<= x"45";
        when x"017A" => data_out<= x"8C";
        when x"017B" => data_out<= x"A9";
        when x"017C" => data_out<= x"42";
        when x"017D" => data_out<= x"A2";
        when x"017E" => data_out<= x"B6";
        when x"017F" => data_out<= x"20";
        when x"0180" => data_out<= x"22";
        when x"0181" => data_out<= x"81";
        when x"0182" => data_out<= x"20";
        when x"0183" => data_out<= x"45";
        when x"0184" => data_out<= x"8C";
        when x"0185" => data_out<= x"A9";
        when x"0186" => data_out<= x"93";
        when x"0187" => data_out<= x"A2";
        when x"0188" => data_out<= x"B3";
        when x"0189" => data_out<= x"20";
        when x"018A" => data_out<= x"22";
        when x"018B" => data_out<= x"81";
        when x"018C" => data_out<= x"20";
        when x"018D" => data_out<= x"45";
        when x"018E" => data_out<= x"8C";
        when x"018F" => data_out<= x"A9";
        when x"0190" => data_out<= x"34";
        when x"0191" => data_out<= x"A2";
        when x"0192" => data_out<= x"B2";
        when x"0193" => data_out<= x"20";
        when x"0194" => data_out<= x"22";
        when x"0195" => data_out<= x"81";
        when x"0196" => data_out<= x"20";
        when x"0197" => data_out<= x"91";
        when x"0198" => data_out<= x"8C";
        when x"0199" => data_out<= x"20";
        when x"019A" => data_out<= x"BB";
        when x"019B" => data_out<= x"9E";
        when x"019C" => data_out<= x"A9";
        when x"019D" => data_out<= x"06";
        when x"019E" => data_out<= x"A2";
        when x"019F" => data_out<= x"02";
        when x"01A0" => data_out<= x"20";
        when x"01A1" => data_out<= x"AE";
        when x"01A2" => data_out<= x"81";
        when x"01A3" => data_out<= x"A0";
        when x"01A4" => data_out<= x"00";
        when x"01A5" => data_out<= x"91";
        when x"01A6" => data_out<= x"0C";
        when x"01A7" => data_out<= x"C9";
        when x"01A8" => data_out<= x"02";
        when x"01A9" => data_out<= x"D0";
        when x"01AA" => data_out<= x"EB";
        when x"01AB" => data_out<= x"4C";
        when x"01AC" => data_out<= x"05";
        when x"01AD" => data_out<= x"AF";
        when x"01AE" => data_out<= x"20";
        when x"01AF" => data_out<= x"7B";
        when x"01B0" => data_out<= x"B0";
        when x"01B1" => data_out<= x"A0";
        when x"01B2" => data_out<= x"16";
        when x"01B3" => data_out<= x"20";
        when x"01B4" => data_out<= x"13";
        when x"01B5" => data_out<= x"B1";
        when x"01B6" => data_out<= x"4C";
        when x"01B7" => data_out<= x"C6";
        when x"01B8" => data_out<= x"81";
        when x"01B9" => data_out<= x"A0";
        when x"01BA" => data_out<= x"17";
        when x"01BB" => data_out<= x"20";
        when x"01BC" => data_out<= x"4F";
        when x"01BD" => data_out<= x"AF";
        when x"01BE" => data_out<= x"20";
        when x"01BF" => data_out<= x"E2";
        when x"01C0" => data_out<= x"AE";
        when x"01C1" => data_out<= x"A0";
        when x"01C2" => data_out<= x"16";
        when x"01C3" => data_out<= x"20";
        when x"01C4" => data_out<= x"C5";
        when x"01C5" => data_out<= x"B0";
        when x"01C6" => data_out<= x"A0";
        when x"01C7" => data_out<= x"17";
        when x"01C8" => data_out<= x"20";
        when x"01C9" => data_out<= x"4F";
        when x"01CA" => data_out<= x"AF";
        when x"01CB" => data_out<= x"85";
        when x"01CC" => data_out<= x"14";
        when x"01CD" => data_out<= x"86";
        when x"01CE" => data_out<= x"15";
        when x"01CF" => data_out<= x"A0";
        when x"01D0" => data_out<= x"00";
        when x"01D1" => data_out<= x"B1";
        when x"01D2" => data_out<= x"14";
        when x"01D3" => data_out<= x"C9";
        when x"01D4" => data_out<= x"20";
        when x"01D5" => data_out<= x"F0";
        when x"01D6" => data_out<= x"E2";
        when x"01D7" => data_out<= x"A0";
        when x"01D8" => data_out<= x"17";
        when x"01D9" => data_out<= x"20";
        when x"01DA" => data_out<= x"4F";
        when x"01DB" => data_out<= x"AF";
        when x"01DC" => data_out<= x"85";
        when x"01DD" => data_out<= x"14";
        when x"01DE" => data_out<= x"86";
        when x"01DF" => data_out<= x"15";
        when x"01E0" => data_out<= x"A0";
        when x"01E1" => data_out<= x"00";
        when x"01E2" => data_out<= x"B1";
        when x"01E3" => data_out<= x"14";
        when x"01E4" => data_out<= x"D0";
        when x"01E5" => data_out<= x"04";
        when x"01E6" => data_out<= x"AA";
        when x"01E7" => data_out<= x"4C";
        when x"01E8" => data_out<= x"44";
        when x"01E9" => data_out<= x"89";
        when x"01EA" => data_out<= x"A0";
        when x"01EB" => data_out<= x"19";
        when x"01EC" => data_out<= x"20";
        when x"01ED" => data_out<= x"93";
        when x"01EE" => data_out<= x"B0";
        when x"01EF" => data_out<= x"A9";
        when x"01F0" => data_out<= x"9A";
        when x"01F1" => data_out<= x"A2";
        when x"01F2" => data_out<= x"BC";
        when x"01F3" => data_out<= x"20";
        when x"01F4" => data_out<= x"F9";
        when x"01F5" => data_out<= x"9A";
        when x"01F6" => data_out<= x"AA";
        when x"01F7" => data_out<= x"F0";
        when x"01F8" => data_out<= x"77";
        when x"01F9" => data_out<= x"A0";
        when x"01FA" => data_out<= x"17";
        when x"01FB" => data_out<= x"20";
        when x"01FC" => data_out<= x"4F";
        when x"01FD" => data_out<= x"AF";
        when x"01FE" => data_out<= x"20";
        when x"01FF" => data_out<= x"FA";
        when x"0200" => data_out<= x"AE";
        when x"0201" => data_out<= x"A0";
        when x"0202" => data_out<= x"13";
        when x"0203" => data_out<= x"20";
        when x"0204" => data_out<= x"C5";
        when x"0205" => data_out<= x"B0";
        when x"0206" => data_out<= x"20";
        when x"0207" => data_out<= x"7B";
        when x"0208" => data_out<= x"B0";
        when x"0209" => data_out<= x"A9";
        when x"020A" => data_out<= x"02";
        when x"020B" => data_out<= x"20";
        when x"020C" => data_out<= x"69";
        when x"020D" => data_out<= x"AF";
        when x"020E" => data_out<= x"20";
        when x"020F" => data_out<= x"7B";
        when x"0210" => data_out<= x"B0";
        when x"0211" => data_out<= x"A9";
        when x"0212" => data_out<= x"0D";
        when x"0213" => data_out<= x"20";
        when x"0214" => data_out<= x"F8";
        when x"0215" => data_out<= x"9D";
        when x"0216" => data_out<= x"A0";
        when x"0217" => data_out<= x"13";
        when x"0218" => data_out<= x"20";
        when x"0219" => data_out<= x"C5";
        when x"021A" => data_out<= x"B0";
        when x"021B" => data_out<= x"20";
        when x"021C" => data_out<= x"7B";
        when x"021D" => data_out<= x"B0";
        when x"021E" => data_out<= x"A9";
        when x"021F" => data_out<= x"13";
        when x"0220" => data_out<= x"20";
        when x"0221" => data_out<= x"69";
        when x"0222" => data_out<= x"AF";
        when x"0223" => data_out<= x"20";
        when x"0224" => data_out<= x"50";
        when x"0225" => data_out<= x"8D";
        when x"0226" => data_out<= x"A0";
        when x"0227" => data_out<= x"13";
        when x"0228" => data_out<= x"20";
        when x"0229" => data_out<= x"C5";
        when x"022A" => data_out<= x"B0";
        when x"022B" => data_out<= x"20";
        when x"022C" => data_out<= x"7B";
        when x"022D" => data_out<= x"B0";
        when x"022E" => data_out<= x"A9";
        when x"022F" => data_out<= x"11";
        when x"0230" => data_out<= x"20";
        when x"0231" => data_out<= x"69";
        when x"0232" => data_out<= x"AF";
        when x"0233" => data_out<= x"20";
        when x"0234" => data_out<= x"50";
        when x"0235" => data_out<= x"8D";
        when x"0236" => data_out<= x"A0";
        when x"0237" => data_out<= x"13";
        when x"0238" => data_out<= x"20";
        when x"0239" => data_out<= x"C5";
        when x"023A" => data_out<= x"B0";
        when x"023B" => data_out<= x"A0";
        when x"023C" => data_out<= x"00";
        when x"023D" => data_out<= x"B1";
        when x"023E" => data_out<= x"0C";
        when x"023F" => data_out<= x"F0";
        when x"0240" => data_out<= x"28";
        when x"0241" => data_out<= x"A0";
        when x"0242" => data_out<= x"12";
        when x"0243" => data_out<= x"B1";
        when x"0244" => data_out<= x"0C";
        when x"0245" => data_out<= x"88";
        when x"0246" => data_out<= x"11";
        when x"0247" => data_out<= x"0C";
        when x"0248" => data_out<= x"F0";
        when x"0249" => data_out<= x"1F";
        when x"024A" => data_out<= x"88";
        when x"024B" => data_out<= x"B1";
        when x"024C" => data_out<= x"0C";
        when x"024D" => data_out<= x"88";
        when x"024E" => data_out<= x"11";
        when x"024F" => data_out<= x"0C";
        when x"0250" => data_out<= x"F0";
        when x"0251" => data_out<= x"17";
        when x"0252" => data_out<= x"A5";
        when x"0253" => data_out<= x"0C";
        when x"0254" => data_out<= x"A6";
        when x"0255" => data_out<= x"0D";
        when x"0256" => data_out<= x"20";
        when x"0257" => data_out<= x"7B";
        when x"0258" => data_out<= x"B0";
        when x"0259" => data_out<= x"A0";
        when x"025A" => data_out<= x"16";
        when x"025B" => data_out<= x"20";
        when x"025C" => data_out<= x"93";
        when x"025D" => data_out<= x"B0";
        when x"025E" => data_out<= x"A0";
        when x"025F" => data_out<= x"14";
        when x"0260" => data_out<= x"20";
        when x"0261" => data_out<= x"4F";
        when x"0262" => data_out<= x"AF";
        when x"0263" => data_out<= x"20";
        when x"0264" => data_out<= x"2B";
        when x"0265" => data_out<= x"96";
        when x"0266" => data_out<= x"4C";
        when x"0267" => data_out<= x"41";
        when x"0268" => data_out<= x"89";
        when x"0269" => data_out<= x"A9";
        when x"026A" => data_out<= x"92";
        when x"026B" => data_out<= x"A2";
        when x"026C" => data_out<= x"B6";
        when x"026D" => data_out<= x"4C";
        when x"026E" => data_out<= x"3E";
        when x"026F" => data_out<= x"89";
        when x"0270" => data_out<= x"A0";
        when x"0271" => data_out<= x"19";
        when x"0272" => data_out<= x"20";
        when x"0273" => data_out<= x"93";
        when x"0274" => data_out<= x"B0";
        when x"0275" => data_out<= x"A9";
        when x"0276" => data_out<= x"95";
        when x"0277" => data_out<= x"A2";
        when x"0278" => data_out<= x"BC";
        when x"0279" => data_out<= x"20";
        when x"027A" => data_out<= x"F9";
        when x"027B" => data_out<= x"9A";
        when x"027C" => data_out<= x"AA";
        when x"027D" => data_out<= x"F0";
        when x"027E" => data_out<= x"60";
        when x"027F" => data_out<= x"A0";
        when x"0280" => data_out<= x"17";
        when x"0281" => data_out<= x"20";
        when x"0282" => data_out<= x"4F";
        when x"0283" => data_out<= x"AF";
        when x"0284" => data_out<= x"20";
        when x"0285" => data_out<= x"FA";
        when x"0286" => data_out<= x"AE";
        when x"0287" => data_out<= x"A0";
        when x"0288" => data_out<= x"13";
        when x"0289" => data_out<= x"20";
        when x"028A" => data_out<= x"C5";
        when x"028B" => data_out<= x"B0";
        when x"028C" => data_out<= x"20";
        when x"028D" => data_out<= x"7B";
        when x"028E" => data_out<= x"B0";
        when x"028F" => data_out<= x"A9";
        when x"0290" => data_out<= x"02";
        when x"0291" => data_out<= x"20";
        when x"0292" => data_out<= x"69";
        when x"0293" => data_out<= x"AF";
        when x"0294" => data_out<= x"20";
        when x"0295" => data_out<= x"7B";
        when x"0296" => data_out<= x"B0";
        when x"0297" => data_out<= x"A9";
        when x"0298" => data_out<= x"0D";
        when x"0299" => data_out<= x"20";
        when x"029A" => data_out<= x"F8";
        when x"029B" => data_out<= x"9D";
        when x"029C" => data_out<= x"A0";
        when x"029D" => data_out<= x"13";
        when x"029E" => data_out<= x"20";
        when x"029F" => data_out<= x"C5";
        when x"02A0" => data_out<= x"B0";
        when x"02A1" => data_out<= x"20";
        when x"02A2" => data_out<= x"7B";
        when x"02A3" => data_out<= x"B0";
        when x"02A4" => data_out<= x"A9";
        when x"02A5" => data_out<= x"13";
        when x"02A6" => data_out<= x"20";
        when x"02A7" => data_out<= x"69";
        when x"02A8" => data_out<= x"AF";
        when x"02A9" => data_out<= x"20";
        when x"02AA" => data_out<= x"50";
        when x"02AB" => data_out<= x"8D";
        when x"02AC" => data_out<= x"A0";
        when x"02AD" => data_out<= x"13";
        when x"02AE" => data_out<= x"20";
        when x"02AF" => data_out<= x"C5";
        when x"02B0" => data_out<= x"B0";
        when x"02B1" => data_out<= x"A0";
        when x"02B2" => data_out<= x"11";
        when x"02B3" => data_out<= x"B1";
        when x"02B4" => data_out<= x"0C";
        when x"02B5" => data_out<= x"C8";
        when x"02B6" => data_out<= x"11";
        when x"02B7" => data_out<= x"0C";
        when x"02B8" => data_out<= x"D0";
        when x"02B9" => data_out<= x"06";
        when x"02BA" => data_out<= x"A2";
        when x"02BB" => data_out<= x"08";
        when x"02BC" => data_out<= x"88";
        when x"02BD" => data_out<= x"20";
        when x"02BE" => data_out<= x"C5";
        when x"02BF" => data_out<= x"B0";
        when x"02C0" => data_out<= x"A0";
        when x"02C1" => data_out<= x"00";
        when x"02C2" => data_out<= x"B1";
        when x"02C3" => data_out<= x"0C";
        when x"02C4" => data_out<= x"F0";
        when x"02C5" => data_out<= x"12";
        when x"02C6" => data_out<= x"A5";
        when x"02C7" => data_out<= x"0C";
        when x"02C8" => data_out<= x"A6";
        when x"02C9" => data_out<= x"0D";
        when x"02CA" => data_out<= x"20";
        when x"02CB" => data_out<= x"7B";
        when x"02CC" => data_out<= x"B0";
        when x"02CD" => data_out<= x"A0";
        when x"02CE" => data_out<= x"14";
        when x"02CF" => data_out<= x"20";
        when x"02D0" => data_out<= x"4F";
        when x"02D1" => data_out<= x"AF";
        when x"02D2" => data_out<= x"20";
        when x"02D3" => data_out<= x"AF";
        when x"02D4" => data_out<= x"97";
        when x"02D5" => data_out<= x"4C";
        when x"02D6" => data_out<= x"41";
        when x"02D7" => data_out<= x"89";
        when x"02D8" => data_out<= x"A9";
        when x"02D9" => data_out<= x"AE";
        when x"02DA" => data_out<= x"A2";
        when x"02DB" => data_out<= x"B7";
        when x"02DC" => data_out<= x"4C";
        when x"02DD" => data_out<= x"3E";
        when x"02DE" => data_out<= x"89";
        when x"02DF" => data_out<= x"A0";
        when x"02E0" => data_out<= x"19";
        when x"02E1" => data_out<= x"20";
        when x"02E2" => data_out<= x"93";
        when x"02E3" => data_out<= x"B0";
        when x"02E4" => data_out<= x"A9";
        when x"02E5" => data_out<= x"11";
        when x"02E6" => data_out<= x"A2";
        when x"02E7" => data_out<= x"BD";
        when x"02E8" => data_out<= x"20";
        when x"02E9" => data_out<= x"F9";
        when x"02EA" => data_out<= x"9A";
        when x"02EB" => data_out<= x"AA";
        when x"02EC" => data_out<= x"F0";
        when x"02ED" => data_out<= x"39";
        when x"02EE" => data_out<= x"A0";
        when x"02EF" => data_out<= x"17";
        when x"02F0" => data_out<= x"20";
        when x"02F1" => data_out<= x"4F";
        when x"02F2" => data_out<= x"AF";
        when x"02F3" => data_out<= x"20";
        when x"02F4" => data_out<= x"F0";
        when x"02F5" => data_out<= x"AE";
        when x"02F6" => data_out<= x"A0";
        when x"02F7" => data_out<= x"13";
        when x"02F8" => data_out<= x"20";
        when x"02F9" => data_out<= x"C5";
        when x"02FA" => data_out<= x"B0";
        when x"02FB" => data_out<= x"20";
        when x"02FC" => data_out<= x"7B";
        when x"02FD" => data_out<= x"B0";
        when x"02FE" => data_out<= x"A9";
        when x"02FF" => data_out<= x"02";
        when x"0300" => data_out<= x"20";
        when x"0301" => data_out<= x"69";
        when x"0302" => data_out<= x"AF";
        when x"0303" => data_out<= x"20";
        when x"0304" => data_out<= x"7B";
        when x"0305" => data_out<= x"B0";
        when x"0306" => data_out<= x"A9";
        when x"0307" => data_out<= x"0D";
        when x"0308" => data_out<= x"20";
        when x"0309" => data_out<= x"F8";
        when x"030A" => data_out<= x"9D";
        when x"030B" => data_out<= x"A0";
        when x"030C" => data_out<= x"13";
        when x"030D" => data_out<= x"20";
        when x"030E" => data_out<= x"C5";
        when x"030F" => data_out<= x"B0";
        when x"0310" => data_out<= x"A0";
        when x"0311" => data_out<= x"00";
        when x"0312" => data_out<= x"B1";
        when x"0313" => data_out<= x"0C";
        when x"0314" => data_out<= x"F0";
        when x"0315" => data_out<= x"0A";
        when x"0316" => data_out<= x"A5";
        when x"0317" => data_out<= x"0C";
        when x"0318" => data_out<= x"A6";
        when x"0319" => data_out<= x"0D";
        when x"031A" => data_out<= x"20";
        when x"031B" => data_out<= x"2A";
        when x"031C" => data_out<= x"99";
        when x"031D" => data_out<= x"4C";
        when x"031E" => data_out<= x"41";
        when x"031F" => data_out<= x"89";
        when x"0320" => data_out<= x"A9";
        when x"0321" => data_out<= x"07";
        when x"0322" => data_out<= x"A2";
        when x"0323" => data_out<= x"BB";
        when x"0324" => data_out<= x"4C";
        when x"0325" => data_out<= x"3E";
        when x"0326" => data_out<= x"89";
        when x"0327" => data_out<= x"A0";
        when x"0328" => data_out<= x"19";
        when x"0329" => data_out<= x"20";
        when x"032A" => data_out<= x"93";
        when x"032B" => data_out<= x"B0";
        when x"032C" => data_out<= x"A9";
        when x"032D" => data_out<= x"39";
        when x"032E" => data_out<= x"A2";
        when x"032F" => data_out<= x"BD";
        when x"0330" => data_out<= x"20";
        when x"0331" => data_out<= x"F9";
        when x"0332" => data_out<= x"9A";
        when x"0333" => data_out<= x"AA";
        when x"0334" => data_out<= x"F0";
        when x"0335" => data_out<= x"39";
        when x"0336" => data_out<= x"A0";
        when x"0337" => data_out<= x"17";
        when x"0338" => data_out<= x"20";
        when x"0339" => data_out<= x"4F";
        when x"033A" => data_out<= x"AF";
        when x"033B" => data_out<= x"20";
        when x"033C" => data_out<= x"F0";
        when x"033D" => data_out<= x"AE";
        when x"033E" => data_out<= x"A0";
        when x"033F" => data_out<= x"13";
        when x"0340" => data_out<= x"20";
        when x"0341" => data_out<= x"C5";
        when x"0342" => data_out<= x"B0";
        when x"0343" => data_out<= x"20";
        when x"0344" => data_out<= x"7B";
        when x"0345" => data_out<= x"B0";
        when x"0346" => data_out<= x"A9";
        when x"0347" => data_out<= x"02";
        when x"0348" => data_out<= x"20";
        when x"0349" => data_out<= x"69";
        when x"034A" => data_out<= x"AF";
        when x"034B" => data_out<= x"20";
        when x"034C" => data_out<= x"7B";
        when x"034D" => data_out<= x"B0";
        when x"034E" => data_out<= x"A9";
        when x"034F" => data_out<= x"0D";
        when x"0350" => data_out<= x"20";
        when x"0351" => data_out<= x"F8";
        when x"0352" => data_out<= x"9D";
        when x"0353" => data_out<= x"A0";
        when x"0354" => data_out<= x"13";
        when x"0355" => data_out<= x"20";
        when x"0356" => data_out<= x"C5";
        when x"0357" => data_out<= x"B0";
        when x"0358" => data_out<= x"A0";
        when x"0359" => data_out<= x"00";
        when x"035A" => data_out<= x"B1";
        when x"035B" => data_out<= x"0C";
        when x"035C" => data_out<= x"F0";
        when x"035D" => data_out<= x"0A";
        when x"035E" => data_out<= x"A5";
        when x"035F" => data_out<= x"0C";
        when x"0360" => data_out<= x"A6";
        when x"0361" => data_out<= x"0D";
        when x"0362" => data_out<= x"20";
        when x"0363" => data_out<= x"75";
        when x"0364" => data_out<= x"99";
        when x"0365" => data_out<= x"4C";
        when x"0366" => data_out<= x"41";
        when x"0367" => data_out<= x"89";
        when x"0368" => data_out<= x"A9";
        when x"0369" => data_out<= x"F7";
        when x"036A" => data_out<= x"A2";
        when x"036B" => data_out<= x"BA";
        when x"036C" => data_out<= x"4C";
        when x"036D" => data_out<= x"3E";
        when x"036E" => data_out<= x"89";
        when x"036F" => data_out<= x"A0";
        when x"0370" => data_out<= x"19";
        when x"0371" => data_out<= x"20";
        when x"0372" => data_out<= x"93";
        when x"0373" => data_out<= x"B0";
        when x"0374" => data_out<= x"A9";
        when x"0375" => data_out<= x"80";
        when x"0376" => data_out<= x"A2";
        when x"0377" => data_out<= x"BD";
        when x"0378" => data_out<= x"20";
        when x"0379" => data_out<= x"F9";
        when x"037A" => data_out<= x"9A";
        when x"037B" => data_out<= x"AA";
        when x"037C" => data_out<= x"F0";
        when x"037D" => data_out<= x"06";
        when x"037E" => data_out<= x"20";
        when x"037F" => data_out<= x"87";
        when x"0380" => data_out<= x"95";
        when x"0381" => data_out<= x"4C";
        when x"0382" => data_out<= x"41";
        when x"0383" => data_out<= x"89";
        when x"0384" => data_out<= x"A0";
        when x"0385" => data_out<= x"19";
        when x"0386" => data_out<= x"20";
        when x"0387" => data_out<= x"93";
        when x"0388" => data_out<= x"B0";
        when x"0389" => data_out<= x"A9";
        when x"038A" => data_out<= x"3F";
        when x"038B" => data_out<= x"A2";
        when x"038C" => data_out<= x"B6";
        when x"038D" => data_out<= x"20";
        when x"038E" => data_out<= x"F9";
        when x"038F" => data_out<= x"9A";
        when x"0390" => data_out<= x"AA";
        when x"0391" => data_out<= x"F0";
        when x"0392" => data_out<= x"06";
        when x"0393" => data_out<= x"20";
        when x"0394" => data_out<= x"B7";
        when x"0395" => data_out<= x"94";
        when x"0396" => data_out<= x"4C";
        when x"0397" => data_out<= x"41";
        when x"0398" => data_out<= x"89";
        when x"0399" => data_out<= x"A0";
        when x"039A" => data_out<= x"19";
        when x"039B" => data_out<= x"20";
        when x"039C" => data_out<= x"93";
        when x"039D" => data_out<= x"B0";
        when x"039E" => data_out<= x"A9";
        when x"039F" => data_out<= x"0A";
        when x"03A0" => data_out<= x"A2";
        when x"03A1" => data_out<= x"BC";
        when x"03A2" => data_out<= x"20";
        when x"03A3" => data_out<= x"F9";
        when x"03A4" => data_out<= x"9A";
        when x"03A5" => data_out<= x"AA";
        when x"03A6" => data_out<= x"F0";
        when x"03A7" => data_out<= x"3C";
        when x"03A8" => data_out<= x"20";
        when x"03A9" => data_out<= x"6A";
        when x"03AA" => data_out<= x"AE";
        when x"03AB" => data_out<= x"A9";
        when x"03AC" => data_out<= x"5E";
        when x"03AD" => data_out<= x"A2";
        when x"03AE" => data_out<= x"BA";
        when x"03AF" => data_out<= x"20";
        when x"03B0" => data_out<= x"22";
        when x"03B1" => data_out<= x"81";
        when x"03B2" => data_out<= x"20";
        when x"03B3" => data_out<= x"45";
        when x"03B4" => data_out<= x"8C";
        when x"03B5" => data_out<= x"20";
        when x"03B6" => data_out<= x"9D";
        when x"03B7" => data_out<= x"A3";
        when x"03B8" => data_out<= x"A0";
        when x"03B9" => data_out<= x"00";
        when x"03BA" => data_out<= x"91";
        when x"03BB" => data_out<= x"0C";
        when x"03BC" => data_out<= x"B1";
        when x"03BD" => data_out<= x"0C";
        when x"03BE" => data_out<= x"D0";
        when x"03BF" => data_out<= x"0A";
        when x"03C0" => data_out<= x"A9";
        when x"03C1" => data_out<= x"94";
        when x"03C2" => data_out<= x"A2";
        when x"03C3" => data_out<= x"BA";
        when x"03C4" => data_out<= x"20";
        when x"03C5" => data_out<= x"22";
        when x"03C6" => data_out<= x"81";
        when x"03C7" => data_out<= x"4C";
        when x"03C8" => data_out<= x"D8";
        when x"03C9" => data_out<= x"83";
        when x"03CA" => data_out<= x"A9";
        when x"03CB" => data_out<= x"2C";
        when x"03CC" => data_out<= x"A2";
        when x"03CD" => data_out<= x"BC";
        when x"03CE" => data_out<= x"20";
        when x"03CF" => data_out<= x"22";
        when x"03D0" => data_out<= x"81";
        when x"03D1" => data_out<= x"A0";
        when x"03D2" => data_out<= x"00";
        when x"03D3" => data_out<= x"B1";
        when x"03D4" => data_out<= x"0C";
        when x"03D5" => data_out<= x"20";
        when x"03D6" => data_out<= x"FD";
        when x"03D7" => data_out<= x"8B";
        when x"03D8" => data_out<= x"20";
        when x"03D9" => data_out<= x"45";
        when x"03DA" => data_out<= x"8C";
        when x"03DB" => data_out<= x"A2";
        when x"03DC" => data_out<= x"00";
        when x"03DD" => data_out<= x"8A";
        when x"03DE" => data_out<= x"20";
        when x"03DF" => data_out<= x"05";
        when x"03E0" => data_out<= x"AF";
        when x"03E1" => data_out<= x"4C";
        when x"03E2" => data_out<= x"44";
        when x"03E3" => data_out<= x"89";
        when x"03E4" => data_out<= x"A0";
        when x"03E5" => data_out<= x"19";
        when x"03E6" => data_out<= x"20";
        when x"03E7" => data_out<= x"93";
        when x"03E8" => data_out<= x"B0";
        when x"03E9" => data_out<= x"A9";
        when x"03EA" => data_out<= x"61";
        when x"03EB" => data_out<= x"A2";
        when x"03EC" => data_out<= x"BC";
        when x"03ED" => data_out<= x"20";
        when x"03EE" => data_out<= x"F9";
        when x"03EF" => data_out<= x"9A";
        when x"03F0" => data_out<= x"AA";
        when x"03F1" => data_out<= x"D0";
        when x"03F2" => data_out<= x"03";
        when x"03F3" => data_out<= x"4C";
        when x"03F4" => data_out<= x"E7";
        when x"03F5" => data_out<= x"84";
        when x"03F6" => data_out<= x"20";
        when x"03F7" => data_out<= x"73";
        when x"03F8" => data_out<= x"AE";
        when x"03F9" => data_out<= x"A0";
        when x"03FA" => data_out<= x"19";
        when x"03FB" => data_out<= x"20";
        when x"03FC" => data_out<= x"4F";
        when x"03FD" => data_out<= x"AF";
        when x"03FE" => data_out<= x"20";
        when x"03FF" => data_out<= x"F5";
        when x"0400" => data_out<= x"AE";
        when x"0401" => data_out<= x"A0";
        when x"0402" => data_out<= x"15";
        when x"0403" => data_out<= x"20";
        when x"0404" => data_out<= x"C5";
        when x"0405" => data_out<= x"B0";
        when x"0406" => data_out<= x"20";
        when x"0407" => data_out<= x"7B";
        when x"0408" => data_out<= x"B0";
        when x"0409" => data_out<= x"A9";
        when x"040A" => data_out<= x"15";
        when x"040B" => data_out<= x"20";
        when x"040C" => data_out<= x"69";
        when x"040D" => data_out<= x"AF";
        when x"040E" => data_out<= x"20";
        when x"040F" => data_out<= x"50";
        when x"0410" => data_out<= x"8D";
        when x"0411" => data_out<= x"A0";
        when x"0412" => data_out<= x"15";
        when x"0413" => data_out<= x"20";
        when x"0414" => data_out<= x"C5";
        when x"0415" => data_out<= x"B0";
        when x"0416" => data_out<= x"A0";
        when x"0417" => data_out<= x"13";
        when x"0418" => data_out<= x"B1";
        when x"0419" => data_out<= x"0C";
        when x"041A" => data_out<= x"C8";
        when x"041B" => data_out<= x"11";
        when x"041C" => data_out<= x"0C";
        when x"041D" => data_out<= x"D0";
        when x"041E" => data_out<= x"06";
        when x"041F" => data_out<= x"A2";
        when x"0420" => data_out<= x"08";
        when x"0421" => data_out<= x"88";
        when x"0422" => data_out<= x"20";
        when x"0423" => data_out<= x"C5";
        when x"0424" => data_out<= x"B0";
        when x"0425" => data_out<= x"A9";
        when x"0426" => data_out<= x"FB";
        when x"0427" => data_out<= x"A2";
        when x"0428" => data_out<= x"B8";
        when x"0429" => data_out<= x"20";
        when x"042A" => data_out<= x"22";
        when x"042B" => data_out<= x"81";
        when x"042C" => data_out<= x"A0";
        when x"042D" => data_out<= x"14";
        when x"042E" => data_out<= x"20";
        when x"042F" => data_out<= x"4F";
        when x"0430" => data_out<= x"AF";
        when x"0431" => data_out<= x"20";
        when x"0432" => data_out<= x"31";
        when x"0433" => data_out<= x"8C";
        when x"0434" => data_out<= x"20";
        when x"0435" => data_out<= x"45";
        when x"0436" => data_out<= x"8C";
        when x"0437" => data_out<= x"A9";
        when x"0438" => data_out<= x"56";
        when x"0439" => data_out<= x"A2";
        when x"043A" => data_out<= x"B8";
        when x"043B" => data_out<= x"20";
        when x"043C" => data_out<= x"22";
        when x"043D" => data_out<= x"81";
        when x"043E" => data_out<= x"20";
        when x"043F" => data_out<= x"45";
        when x"0440" => data_out<= x"8C";
        when x"0441" => data_out<= x"A0";
        when x"0442" => data_out<= x"14";
        when x"0443" => data_out<= x"20";
        when x"0444" => data_out<= x"4F";
        when x"0445" => data_out<= x"AF";
        when x"0446" => data_out<= x"20";
        when x"0447" => data_out<= x"C7";
        when x"0448" => data_out<= x"AB";
        when x"0449" => data_out<= x"20";
        when x"044A" => data_out<= x"C3";
        when x"044B" => data_out<= x"B0";
        when x"044C" => data_out<= x"20";
        when x"044D" => data_out<= x"73";
        when x"044E" => data_out<= x"AE";
        when x"044F" => data_out<= x"A2";
        when x"0450" => data_out<= x"00";
        when x"0451" => data_out<= x"8A";
        when x"0452" => data_out<= x"20";
        when x"0453" => data_out<= x"C3";
        when x"0454" => data_out<= x"B0";
        when x"0455" => data_out<= x"A0";
        when x"0456" => data_out<= x"01";
        when x"0457" => data_out<= x"B1";
        when x"0458" => data_out<= x"0C";
        when x"0459" => data_out<= x"C9";
        when x"045A" => data_out<= x"75";
        when x"045B" => data_out<= x"D0";
        when x"045C" => data_out<= x"05";
        when x"045D" => data_out<= x"88";
        when x"045E" => data_out<= x"B1";
        when x"045F" => data_out<= x"0C";
        when x"0460" => data_out<= x"C9";
        when x"0461" => data_out<= x"30";
        when x"0462" => data_out<= x"B0";
        when x"0463" => data_out<= x"09";
        when x"0464" => data_out<= x"20";
        when x"0465" => data_out<= x"4D";
        when x"0466" => data_out<= x"AF";
        when x"0467" => data_out<= x"20";
        when x"0468" => data_out<= x"E2";
        when x"0469" => data_out<= x"AE";
        when x"046A" => data_out<= x"4C";
        when x"046B" => data_out<= x"52";
        when x"046C" => data_out<= x"84";
        when x"046D" => data_out<= x"20";
        when x"046E" => data_out<= x"14";
        when x"046F" => data_out<= x"AF";
        when x"0470" => data_out<= x"4C";
        when x"0471" => data_out<= x"76";
        when x"0472" => data_out<= x"84";
        when x"0473" => data_out<= x"20";
        when x"0474" => data_out<= x"FD";
        when x"0475" => data_out<= x"80";
        when x"0476" => data_out<= x"20";
        when x"0477" => data_out<= x"0A";
        when x"0478" => data_out<= x"81";
        when x"0479" => data_out<= x"AA";
        when x"047A" => data_out<= x"D0";
        when x"047B" => data_out<= x"F7";
        when x"047C" => data_out<= x"20";
        when x"047D" => data_out<= x"4D";
        when x"047E" => data_out<= x"AF";
        when x"047F" => data_out<= x"C9";
        when x"0480" => data_out<= x"01";
        when x"0481" => data_out<= x"8A";
        when x"0482" => data_out<= x"E9";
        when x"0483" => data_out<= x"00";
        when x"0484" => data_out<= x"70";
        when x"0485" => data_out<= x"02";
        when x"0486" => data_out<= x"49";
        when x"0487" => data_out<= x"80";
        when x"0488" => data_out<= x"10";
        when x"0489" => data_out<= x"3E";
        when x"048A" => data_out<= x"20";
        when x"048B" => data_out<= x"45";
        when x"048C" => data_out<= x"8C";
        when x"048D" => data_out<= x"A9";
        when x"048E" => data_out<= x"A4";
        when x"048F" => data_out<= x"A2";
        when x"0490" => data_out<= x"BC";
        when x"0491" => data_out<= x"20";
        when x"0492" => data_out<= x"22";
        when x"0493" => data_out<= x"81";
        when x"0494" => data_out<= x"20";
        when x"0495" => data_out<= x"4D";
        when x"0496" => data_out<= x"AF";
        when x"0497" => data_out<= x"20";
        when x"0498" => data_out<= x"86";
        when x"0499" => data_out<= x"93";
        when x"049A" => data_out<= x"A9";
        when x"049B" => data_out<= x"CA";
        when x"049C" => data_out<= x"A2";
        when x"049D" => data_out<= x"BB";
        when x"049E" => data_out<= x"20";
        when x"049F" => data_out<= x"22";
        when x"04A0" => data_out<= x"81";
        when x"04A1" => data_out<= x"A0";
        when x"04A2" => data_out<= x"14";
        when x"04A3" => data_out<= x"20";
        when x"04A4" => data_out<= x"4F";
        when x"04A5" => data_out<= x"AF";
        when x"04A6" => data_out<= x"20";
        when x"04A7" => data_out<= x"31";
        when x"04A8" => data_out<= x"8C";
        when x"04A9" => data_out<= x"A9";
        when x"04AA" => data_out<= x"7D";
        when x"04AB" => data_out<= x"A2";
        when x"04AC" => data_out<= x"BD";
        when x"04AD" => data_out<= x"20";
        when x"04AE" => data_out<= x"22";
        when x"04AF" => data_out<= x"81";
        when x"04B0" => data_out<= x"20";
        when x"04B1" => data_out<= x"4D";
        when x"04B2" => data_out<= x"AF";
        when x"04B3" => data_out<= x"18";
        when x"04B4" => data_out<= x"A0";
        when x"04B5" => data_out<= x"13";
        when x"04B6" => data_out<= x"71";
        when x"04B7" => data_out<= x"0C";
        when x"04B8" => data_out<= x"48";
        when x"04B9" => data_out<= x"8A";
        when x"04BA" => data_out<= x"C8";
        when x"04BB" => data_out<= x"71";
        when x"04BC" => data_out<= x"0C";
        when x"04BD" => data_out<= x"AA";
        when x"04BE" => data_out<= x"68";
        when x"04BF" => data_out<= x"20";
        when x"04C0" => data_out<= x"5A";
        when x"04C1" => data_out<= x"AE";
        when x"04C2" => data_out<= x"20";
        when x"04C3" => data_out<= x"31";
        when x"04C4" => data_out<= x"8C";
        when x"04C5" => data_out<= x"4C";
        when x"04C6" => data_out<= x"DB";
        when x"04C7" => data_out<= x"84";
        when x"04C8" => data_out<= x"20";
        when x"04C9" => data_out<= x"45";
        when x"04CA" => data_out<= x"8C";
        when x"04CB" => data_out<= x"A9";
        when x"04CC" => data_out<= x"37";
        when x"04CD" => data_out<= x"A2";
        when x"04CE" => data_out<= x"BB";
        when x"04CF" => data_out<= x"20";
        when x"04D0" => data_out<= x"22";
        when x"04D1" => data_out<= x"81";
        when x"04D2" => data_out<= x"20";
        when x"04D3" => data_out<= x"4D";
        when x"04D4" => data_out<= x"AF";
        when x"04D5" => data_out<= x"20";
        when x"04D6" => data_out<= x"33";
        when x"04D7" => data_out<= x"B0";
        when x"04D8" => data_out<= x"20";
        when x"04D9" => data_out<= x"FD";
        when x"04DA" => data_out<= x"8B";
        when x"04DB" => data_out<= x"20";
        when x"04DC" => data_out<= x"45";
        when x"04DD" => data_out<= x"8C";
        when x"04DE" => data_out<= x"A2";
        when x"04DF" => data_out<= x"00";
        when x"04E0" => data_out<= x"8A";
        when x"04E1" => data_out<= x"20";
        when x"04E2" => data_out<= x"14";
        when x"04E3" => data_out<= x"AF";
        when x"04E4" => data_out<= x"4C";
        when x"04E5" => data_out<= x"44";
        when x"04E6" => data_out<= x"89";
        when x"04E7" => data_out<= x"A0";
        when x"04E8" => data_out<= x"17";
        when x"04E9" => data_out<= x"20";
        when x"04EA" => data_out<= x"4F";
        when x"04EB" => data_out<= x"AF";
        when x"04EC" => data_out<= x"85";
        when x"04ED" => data_out<= x"14";
        when x"04EE" => data_out<= x"86";
        when x"04EF" => data_out<= x"15";
        when x"04F0" => data_out<= x"A0";
        when x"04F1" => data_out<= x"00";
        when x"04F2" => data_out<= x"B1";
        when x"04F3" => data_out<= x"14";
        when x"04F4" => data_out<= x"A0";
        when x"04F5" => data_out<= x"15";
        when x"04F6" => data_out<= x"91";
        when x"04F7" => data_out<= x"0C";
        when x"04F8" => data_out<= x"C9";
        when x"04F9" => data_out<= x"61";
        when x"04FA" => data_out<= x"90";
        when x"04FB" => data_out<= x"0B";
        when x"04FC" => data_out<= x"B1";
        when x"04FD" => data_out<= x"0C";
        when x"04FE" => data_out<= x"C9";
        when x"04FF" => data_out<= x"7B";
        when x"0500" => data_out<= x"B0";
        when x"0501" => data_out<= x"05";
        when x"0502" => data_out<= x"38";
        when x"0503" => data_out<= x"E9";
        when x"0504" => data_out<= x"20";
        when x"0505" => data_out<= x"91";
        when x"0506" => data_out<= x"0C";
        when x"0507" => data_out<= x"A0";
        when x"0508" => data_out<= x"17";
        when x"0509" => data_out<= x"20";
        when x"050A" => data_out<= x"4F";
        when x"050B" => data_out<= x"AF";
        when x"050C" => data_out<= x"20";
        when x"050D" => data_out<= x"E2";
        when x"050E" => data_out<= x"AE";
        when x"050F" => data_out<= x"A0";
        when x"0510" => data_out<= x"13";
        when x"0511" => data_out<= x"20";
        when x"0512" => data_out<= x"C5";
        when x"0513" => data_out<= x"B0";
        when x"0514" => data_out<= x"A0";
        when x"0515" => data_out<= x"15";
        when x"0516" => data_out<= x"B1";
        when x"0517" => data_out<= x"0C";
        when x"0518" => data_out<= x"C9";
        when x"0519" => data_out<= x"3F";
        when x"051A" => data_out<= x"D0";
        when x"051B" => data_out<= x"03";
        when x"051C" => data_out<= x"4C";
        when x"051D" => data_out<= x"9C";
        when x"051E" => data_out<= x"88";
        when x"051F" => data_out<= x"C9";
        when x"0520" => data_out<= x"44";
        when x"0521" => data_out<= x"D0";
        when x"0522" => data_out<= x"03";
        when x"0523" => data_out<= x"4C";
        when x"0524" => data_out<= x"09";
        when x"0525" => data_out<= x"87";
        when x"0526" => data_out<= x"C9";
        when x"0527" => data_out<= x"46";
        when x"0528" => data_out<= x"D0";
        when x"0529" => data_out<= x"03";
        when x"052A" => data_out<= x"4C";
        when x"052B" => data_out<= x"79";
        when x"052C" => data_out<= x"87";
        when x"052D" => data_out<= x"C9";
        when x"052E" => data_out<= x"48";
        when x"052F" => data_out<= x"D0";
        when x"0530" => data_out<= x"03";
        when x"0531" => data_out<= x"4C";
        when x"0532" => data_out<= x"9C";
        when x"0533" => data_out<= x"88";
        when x"0534" => data_out<= x"C9";
        when x"0535" => data_out<= x"49";
        when x"0536" => data_out<= x"D0";
        when x"0537" => data_out<= x"03";
        when x"0538" => data_out<= x"4C";
        when x"0539" => data_out<= x"6E";
        when x"053A" => data_out<= x"88";
        when x"053B" => data_out<= x"C9";
        when x"053C" => data_out<= x"4C";
        when x"053D" => data_out<= x"D0";
        when x"053E" => data_out<= x"03";
        when x"053F" => data_out<= x"4C";
        when x"0540" => data_out<= x"4A";
        when x"0541" => data_out<= x"87";
        when x"0542" => data_out<= x"C9";
        when x"0543" => data_out<= x"4D";
        when x"0544" => data_out<= x"D0";
        when x"0545" => data_out<= x"03";
        when x"0546" => data_out<= x"4C";
        when x"0547" => data_out<= x"FC";
        when x"0548" => data_out<= x"87";
        when x"0549" => data_out<= x"C9";
        when x"054A" => data_out<= x"51";
        when x"054B" => data_out<= x"D0";
        when x"054C" => data_out<= x"03";
        when x"054D" => data_out<= x"4C";
        when x"054E" => data_out<= x"7E";
        when x"054F" => data_out<= x"88";
        when x"0550" => data_out<= x"C9";
        when x"0551" => data_out<= x"52";
        when x"0552" => data_out<= x"F0";
        when x"0553" => data_out<= x"1F";
        when x"0554" => data_out<= x"C9";
        when x"0555" => data_out<= x"53";
        when x"0556" => data_out<= x"D0";
        when x"0557" => data_out<= x"03";
        when x"0558" => data_out<= x"4C";
        when x"0559" => data_out<= x"74";
        when x"055A" => data_out<= x"88";
        when x"055B" => data_out<= x"C9";
        when x"055C" => data_out<= x"54";
        when x"055D" => data_out<= x"D0";
        when x"055E" => data_out<= x"03";
        when x"055F" => data_out<= x"4C";
        when x"0560" => data_out<= x"74";
        when x"0561" => data_out<= x"88";
        when x"0562" => data_out<= x"C9";
        when x"0563" => data_out<= x"56";
        when x"0564" => data_out<= x"D0";
        when x"0565" => data_out<= x"03";
        when x"0566" => data_out<= x"4C";
        when x"0567" => data_out<= x"74";
        when x"0568" => data_out<= x"88";
        when x"0569" => data_out<= x"C9";
        when x"056A" => data_out<= x"57";
        when x"056B" => data_out<= x"D0";
        when x"056C" => data_out<= x"03";
        when x"056D" => data_out<= x"4C";
        when x"056E" => data_out<= x"AD";
        when x"056F" => data_out<= x"86";
        when x"0570" => data_out<= x"4C";
        when x"0571" => data_out<= x"3A";
        when x"0572" => data_out<= x"89";
        when x"0573" => data_out<= x"88";
        when x"0574" => data_out<= x"20";
        when x"0575" => data_out<= x"4F";
        when x"0576" => data_out<= x"AF";
        when x"0577" => data_out<= x"85";
        when x"0578" => data_out<= x"14";
        when x"0579" => data_out<= x"86";
        when x"057A" => data_out<= x"15";
        when x"057B" => data_out<= x"A0";
        when x"057C" => data_out<= x"00";
        when x"057D" => data_out<= x"B1";
        when x"057E" => data_out<= x"14";
        when x"057F" => data_out<= x"C9";
        when x"0580" => data_out<= x"20";
        when x"0581" => data_out<= x"F0";
        when x"0582" => data_out<= x"0F";
        when x"0583" => data_out<= x"A0";
        when x"0584" => data_out<= x"14";
        when x"0585" => data_out<= x"20";
        when x"0586" => data_out<= x"4F";
        when x"0587" => data_out<= x"AF";
        when x"0588" => data_out<= x"85";
        when x"0589" => data_out<= x"14";
        when x"058A" => data_out<= x"86";
        when x"058B" => data_out<= x"15";
        when x"058C" => data_out<= x"A0";
        when x"058D" => data_out<= x"00";
        when x"058E" => data_out<= x"B1";
        when x"058F" => data_out<= x"14";
        when x"0590" => data_out<= x"D0";
        when x"0591" => data_out<= x"27";
        when x"0592" => data_out<= x"A0";
        when x"0593" => data_out<= x"16";
        when x"0594" => data_out<= x"20";
        when x"0595" => data_out<= x"93";
        when x"0596" => data_out<= x"B0";
        when x"0597" => data_out<= x"A9";
        when x"0598" => data_out<= x"13";
        when x"0599" => data_out<= x"20";
        when x"059A" => data_out<= x"69";
        when x"059B" => data_out<= x"AF";
        when x"059C" => data_out<= x"20";
        when x"059D" => data_out<= x"50";
        when x"059E" => data_out<= x"8D";
        when x"059F" => data_out<= x"A0";
        when x"05A0" => data_out<= x"11";
        when x"05A1" => data_out<= x"B1";
        when x"05A2" => data_out<= x"0C";
        when x"05A3" => data_out<= x"C8";
        when x"05A4" => data_out<= x"11";
        when x"05A5" => data_out<= x"0C";
        when x"05A6" => data_out<= x"D0";
        when x"05A7" => data_out<= x"08";
        when x"05A8" => data_out<= x"A2";
        when x"05A9" => data_out<= x"08";
        when x"05AA" => data_out<= x"88";
        when x"05AB" => data_out<= x"20";
        when x"05AC" => data_out<= x"C5";
        when x"05AD" => data_out<= x"B0";
        when x"05AE" => data_out<= x"A0";
        when x"05AF" => data_out<= x"12";
        when x"05B0" => data_out<= x"20";
        when x"05B1" => data_out<= x"4F";
        when x"05B2" => data_out<= x"AF";
        when x"05B3" => data_out<= x"20";
        when x"05B4" => data_out<= x"4F";
        when x"05B5" => data_out<= x"8C";
        when x"05B6" => data_out<= x"4C";
        when x"05B7" => data_out<= x"41";
        when x"05B8" => data_out<= x"89";
        when x"05B9" => data_out<= x"A0";
        when x"05BA" => data_out<= x"14";
        when x"05BB" => data_out<= x"20";
        when x"05BC" => data_out<= x"4F";
        when x"05BD" => data_out<= x"AF";
        when x"05BE" => data_out<= x"85";
        when x"05BF" => data_out<= x"14";
        when x"05C0" => data_out<= x"86";
        when x"05C1" => data_out<= x"15";
        when x"05C2" => data_out<= x"A0";
        when x"05C3" => data_out<= x"00";
        when x"05C4" => data_out<= x"B1";
        when x"05C5" => data_out<= x"14";
        when x"05C6" => data_out<= x"C9";
        when x"05C7" => data_out<= x"44";
        when x"05C8" => data_out<= x"F0";
        when x"05C9" => data_out<= x"14";
        when x"05CA" => data_out<= x"A0";
        when x"05CB" => data_out<= x"14";
        when x"05CC" => data_out<= x"20";
        when x"05CD" => data_out<= x"4F";
        when x"05CE" => data_out<= x"AF";
        when x"05CF" => data_out<= x"85";
        when x"05D0" => data_out<= x"14";
        when x"05D1" => data_out<= x"86";
        when x"05D2" => data_out<= x"15";
        when x"05D3" => data_out<= x"A0";
        when x"05D4" => data_out<= x"00";
        when x"05D5" => data_out<= x"B1";
        when x"05D6" => data_out<= x"14";
        when x"05D7" => data_out<= x"C9";
        when x"05D8" => data_out<= x"64";
        when x"05D9" => data_out<= x"F0";
        when x"05DA" => data_out<= x"03";
        when x"05DB" => data_out<= x"4C";
        when x"05DC" => data_out<= x"81";
        when x"05DD" => data_out<= x"86";
        when x"05DE" => data_out<= x"A0";
        when x"05DF" => data_out<= x"14";
        when x"05E0" => data_out<= x"20";
        when x"05E1" => data_out<= x"4F";
        when x"05E2" => data_out<= x"AF";
        when x"05E3" => data_out<= x"20";
        when x"05E4" => data_out<= x"E2";
        when x"05E5" => data_out<= x"AE";
        when x"05E6" => data_out<= x"85";
        when x"05E7" => data_out<= x"14";
        when x"05E8" => data_out<= x"86";
        when x"05E9" => data_out<= x"15";
        when x"05EA" => data_out<= x"A0";
        when x"05EB" => data_out<= x"00";
        when x"05EC" => data_out<= x"B1";
        when x"05ED" => data_out<= x"14";
        when x"05EE" => data_out<= x"C9";
        when x"05EF" => data_out<= x"20";
        when x"05F0" => data_out<= x"F0";
        when x"05F1" => data_out<= x"12";
        when x"05F2" => data_out<= x"A0";
        when x"05F3" => data_out<= x"14";
        when x"05F4" => data_out<= x"20";
        when x"05F5" => data_out<= x"4F";
        when x"05F6" => data_out<= x"AF";
        when x"05F7" => data_out<= x"20";
        when x"05F8" => data_out<= x"E2";
        when x"05F9" => data_out<= x"AE";
        when x"05FA" => data_out<= x"85";
        when x"05FB" => data_out<= x"14";
        when x"05FC" => data_out<= x"86";
        when x"05FD" => data_out<= x"15";
        when x"05FE" => data_out<= x"A0";
        when x"05FF" => data_out<= x"00";
        when x"0600" => data_out<= x"B1";
        when x"0601" => data_out<= x"14";
        when x"0602" => data_out<= x"D0";
        when x"0603" => data_out<= x"7D";
        when x"0604" => data_out<= x"A0";
        when x"0605" => data_out<= x"14";
        when x"0606" => data_out<= x"20";
        when x"0607" => data_out<= x"4F";
        when x"0608" => data_out<= x"AF";
        when x"0609" => data_out<= x"20";
        when x"060A" => data_out<= x"E2";
        when x"060B" => data_out<= x"AE";
        when x"060C" => data_out<= x"A0";
        when x"060D" => data_out<= x"13";
        when x"060E" => data_out<= x"20";
        when x"060F" => data_out<= x"C5";
        when x"0610" => data_out<= x"B0";
        when x"0611" => data_out<= x"20";
        when x"0612" => data_out<= x"7B";
        when x"0613" => data_out<= x"B0";
        when x"0614" => data_out<= x"A9";
        when x"0615" => data_out<= x"13";
        when x"0616" => data_out<= x"20";
        when x"0617" => data_out<= x"69";
        when x"0618" => data_out<= x"AF";
        when x"0619" => data_out<= x"20";
        when x"061A" => data_out<= x"50";
        when x"061B" => data_out<= x"8D";
        when x"061C" => data_out<= x"A0";
        when x"061D" => data_out<= x"13";
        when x"061E" => data_out<= x"20";
        when x"061F" => data_out<= x"C5";
        when x"0620" => data_out<= x"B0";
        when x"0621" => data_out<= x"A0";
        when x"0622" => data_out<= x"11";
        when x"0623" => data_out<= x"B1";
        when x"0624" => data_out<= x"0C";
        when x"0625" => data_out<= x"C8";
        when x"0626" => data_out<= x"11";
        when x"0627" => data_out<= x"0C";
        when x"0628" => data_out<= x"D0";
        when x"0629" => data_out<= x"24";
        when x"062A" => data_out<= x"A0";
        when x"062B" => data_out<= x"14";
        when x"062C" => data_out<= x"20";
        when x"062D" => data_out<= x"4F";
        when x"062E" => data_out<= x"AF";
        when x"062F" => data_out<= x"85";
        when x"0630" => data_out<= x"14";
        when x"0631" => data_out<= x"86";
        when x"0632" => data_out<= x"15";
        when x"0633" => data_out<= x"A0";
        when x"0634" => data_out<= x"17";
        when x"0635" => data_out<= x"20";
        when x"0636" => data_out<= x"4F";
        when x"0637" => data_out<= x"AF";
        when x"0638" => data_out<= x"20";
        when x"0639" => data_out<= x"E9";
        when x"063A" => data_out<= x"AE";
        when x"063B" => data_out<= x"E4";
        when x"063C" => data_out<= x"15";
        when x"063D" => data_out<= x"D0";
        when x"063E" => data_out<= x"0F";
        when x"063F" => data_out<= x"C5";
        when x"0640" => data_out<= x"14";
        when x"0641" => data_out<= x"D0";
        when x"0642" => data_out<= x"0B";
        when x"0643" => data_out<= x"AD";
        when x"0644" => data_out<= x"00";
        when x"0645" => data_out<= x"02";
        when x"0646" => data_out<= x"AE";
        when x"0647" => data_out<= x"01";
        when x"0648" => data_out<= x"02";
        when x"0649" => data_out<= x"A0";
        when x"064A" => data_out<= x"11";
        when x"064B" => data_out<= x"20";
        when x"064C" => data_out<= x"C5";
        when x"064D" => data_out<= x"B0";
        when x"064E" => data_out<= x"A9";
        when x"064F" => data_out<= x"24";
        when x"0650" => data_out<= x"20";
        when x"0651" => data_out<= x"F0";
        when x"0652" => data_out<= x"80";
        when x"0653" => data_out<= x"A0";
        when x"0654" => data_out<= x"12";
        when x"0655" => data_out<= x"20";
        when x"0656" => data_out<= x"4F";
        when x"0657" => data_out<= x"AF";
        when x"0658" => data_out<= x"20";
        when x"0659" => data_out<= x"31";
        when x"065A" => data_out<= x"8C";
        when x"065B" => data_out<= x"A9";
        when x"065C" => data_out<= x"9F";
        when x"065D" => data_out<= x"A2";
        when x"065E" => data_out<= x"BC";
        when x"065F" => data_out<= x"20";
        when x"0660" => data_out<= x"22";
        when x"0661" => data_out<= x"81";
        when x"0662" => data_out<= x"A0";
        when x"0663" => data_out<= x"12";
        when x"0664" => data_out<= x"20";
        when x"0665" => data_out<= x"4F";
        when x"0666" => data_out<= x"AF";
        when x"0667" => data_out<= x"20";
        when x"0668" => data_out<= x"49";
        when x"0669" => data_out<= x"89";
        when x"066A" => data_out<= x"20";
        when x"066B" => data_out<= x"FD";
        when x"066C" => data_out<= x"8B";
        when x"066D" => data_out<= x"20";
        when x"066E" => data_out<= x"45";
        when x"066F" => data_out<= x"8C";
        when x"0670" => data_out<= x"A0";
        when x"0671" => data_out<= x"12";
        when x"0672" => data_out<= x"20";
        when x"0673" => data_out<= x"4F";
        when x"0674" => data_out<= x"AF";
        when x"0675" => data_out<= x"20";
        when x"0676" => data_out<= x"E2";
        when x"0677" => data_out<= x"AE";
        when x"0678" => data_out<= x"8D";
        when x"0679" => data_out<= x"00";
        when x"067A" => data_out<= x"02";
        when x"067B" => data_out<= x"8E";
        when x"067C" => data_out<= x"01";
        when x"067D" => data_out<= x"02";
        when x"067E" => data_out<= x"4C";
        when x"067F" => data_out<= x"41";
        when x"0680" => data_out<= x"89";
        when x"0681" => data_out<= x"A0";
        when x"0682" => data_out<= x"16";
        when x"0683" => data_out<= x"20";
        when x"0684" => data_out<= x"93";
        when x"0685" => data_out<= x"B0";
        when x"0686" => data_out<= x"A9";
        when x"0687" => data_out<= x"13";
        when x"0688" => data_out<= x"20";
        when x"0689" => data_out<= x"69";
        when x"068A" => data_out<= x"AF";
        when x"068B" => data_out<= x"20";
        when x"068C" => data_out<= x"50";
        when x"068D" => data_out<= x"8D";
        when x"068E" => data_out<= x"A0";
        when x"068F" => data_out<= x"13";
        when x"0690" => data_out<= x"20";
        when x"0691" => data_out<= x"C5";
        when x"0692" => data_out<= x"B0";
        when x"0693" => data_out<= x"A0";
        when x"0694" => data_out<= x"11";
        when x"0695" => data_out<= x"B1";
        when x"0696" => data_out<= x"0C";
        when x"0697" => data_out<= x"C8";
        when x"0698" => data_out<= x"11";
        when x"0699" => data_out<= x"0C";
        when x"069A" => data_out<= x"D0";
        when x"069B" => data_out<= x"08";
        when x"069C" => data_out<= x"A2";
        when x"069D" => data_out<= x"08";
        when x"069E" => data_out<= x"88";
        when x"069F" => data_out<= x"20";
        when x"06A0" => data_out<= x"C5";
        when x"06A1" => data_out<= x"B0";
        when x"06A2" => data_out<= x"A0";
        when x"06A3" => data_out<= x"12";
        when x"06A4" => data_out<= x"20";
        when x"06A5" => data_out<= x"4F";
        when x"06A6" => data_out<= x"AF";
        when x"06A7" => data_out<= x"20";
        when x"06A8" => data_out<= x"4F";
        when x"06A9" => data_out<= x"8C";
        when x"06AA" => data_out<= x"4C";
        when x"06AB" => data_out<= x"41";
        when x"06AC" => data_out<= x"89";
        when x"06AD" => data_out<= x"C8";
        when x"06AE" => data_out<= x"20";
        when x"06AF" => data_out<= x"93";
        when x"06B0" => data_out<= x"B0";
        when x"06B1" => data_out<= x"A9";
        when x"06B2" => data_out<= x"13";
        when x"06B3" => data_out<= x"20";
        when x"06B4" => data_out<= x"69";
        when x"06B5" => data_out<= x"AF";
        when x"06B6" => data_out<= x"20";
        when x"06B7" => data_out<= x"50";
        when x"06B8" => data_out<= x"8D";
        when x"06B9" => data_out<= x"A0";
        when x"06BA" => data_out<= x"13";
        when x"06BB" => data_out<= x"20";
        when x"06BC" => data_out<= x"C5";
        when x"06BD" => data_out<= x"B0";
        when x"06BE" => data_out<= x"20";
        when x"06BF" => data_out<= x"7B";
        when x"06C0" => data_out<= x"B0";
        when x"06C1" => data_out<= x"A9";
        when x"06C2" => data_out<= x"0F";
        when x"06C3" => data_out<= x"20";
        when x"06C4" => data_out<= x"69";
        when x"06C5" => data_out<= x"AF";
        when x"06C6" => data_out<= x"20";
        when x"06C7" => data_out<= x"50";
        when x"06C8" => data_out<= x"8D";
        when x"06C9" => data_out<= x"A0";
        when x"06CA" => data_out<= x"13";
        when x"06CB" => data_out<= x"20";
        when x"06CC" => data_out<= x"C5";
        when x"06CD" => data_out<= x"B0";
        when x"06CE" => data_out<= x"A0";
        when x"06CF" => data_out<= x"14";
        when x"06D0" => data_out<= x"20";
        when x"06D1" => data_out<= x"93";
        when x"06D2" => data_out<= x"B0";
        when x"06D3" => data_out<= x"A0";
        when x"06D4" => data_out<= x"0F";
        when x"06D5" => data_out<= x"B1";
        when x"06D6" => data_out<= x"0C";
        when x"06D7" => data_out<= x"20";
        when x"06D8" => data_out<= x"5A";
        when x"06D9" => data_out<= x"89";
        when x"06DA" => data_out<= x"A9";
        when x"06DB" => data_out<= x"24";
        when x"06DC" => data_out<= x"20";
        when x"06DD" => data_out<= x"F0";
        when x"06DE" => data_out<= x"80";
        when x"06DF" => data_out<= x"A0";
        when x"06E0" => data_out<= x"12";
        when x"06E1" => data_out<= x"20";
        when x"06E2" => data_out<= x"4F";
        when x"06E3" => data_out<= x"AF";
        when x"06E4" => data_out<= x"20";
        when x"06E5" => data_out<= x"31";
        when x"06E6" => data_out<= x"8C";
        when x"06E7" => data_out<= x"A9";
        when x"06E8" => data_out<= x"55";
        when x"06E9" => data_out<= x"A2";
        when x"06EA" => data_out<= x"BC";
        when x"06EB" => data_out<= x"20";
        when x"06EC" => data_out<= x"22";
        when x"06ED" => data_out<= x"81";
        when x"06EE" => data_out<= x"A0";
        when x"06EF" => data_out<= x"0D";
        when x"06F0" => data_out<= x"B1";
        when x"06F1" => data_out<= x"0C";
        when x"06F2" => data_out<= x"20";
        when x"06F3" => data_out<= x"FD";
        when x"06F4" => data_out<= x"8B";
        when x"06F5" => data_out<= x"20";
        when x"06F6" => data_out<= x"45";
        when x"06F7" => data_out<= x"8C";
        when x"06F8" => data_out<= x"A0";
        when x"06F9" => data_out<= x"12";
        when x"06FA" => data_out<= x"20";
        when x"06FB" => data_out<= x"4F";
        when x"06FC" => data_out<= x"AF";
        when x"06FD" => data_out<= x"20";
        when x"06FE" => data_out<= x"E2";
        when x"06FF" => data_out<= x"AE";
        when x"0700" => data_out<= x"8D";
        when x"0701" => data_out<= x"00";
        when x"0702" => data_out<= x"02";
        when x"0703" => data_out<= x"8E";
        when x"0704" => data_out<= x"01";
        when x"0705" => data_out<= x"02";
        when x"0706" => data_out<= x"4C";
        when x"0707" => data_out<= x"41";
        when x"0708" => data_out<= x"89";
        when x"0709" => data_out<= x"C8";
        when x"070A" => data_out<= x"20";
        when x"070B" => data_out<= x"93";
        when x"070C" => data_out<= x"B0";
        when x"070D" => data_out<= x"A9";
        when x"070E" => data_out<= x"13";
        when x"070F" => data_out<= x"20";
        when x"0710" => data_out<= x"69";
        when x"0711" => data_out<= x"AF";
        when x"0712" => data_out<= x"20";
        when x"0713" => data_out<= x"50";
        when x"0714" => data_out<= x"8D";
        when x"0715" => data_out<= x"A0";
        when x"0716" => data_out<= x"13";
        when x"0717" => data_out<= x"20";
        when x"0718" => data_out<= x"C5";
        when x"0719" => data_out<= x"B0";
        when x"071A" => data_out<= x"20";
        when x"071B" => data_out<= x"7B";
        when x"071C" => data_out<= x"B0";
        when x"071D" => data_out<= x"A9";
        when x"071E" => data_out<= x"11";
        when x"071F" => data_out<= x"20";
        when x"0720" => data_out<= x"69";
        when x"0721" => data_out<= x"AF";
        when x"0722" => data_out<= x"20";
        when x"0723" => data_out<= x"50";
        when x"0724" => data_out<= x"8D";
        when x"0725" => data_out<= x"A0";
        when x"0726" => data_out<= x"13";
        when x"0727" => data_out<= x"20";
        when x"0728" => data_out<= x"C5";
        when x"0729" => data_out<= x"B0";
        when x"072A" => data_out<= x"A0";
        when x"072B" => data_out<= x"0F";
        when x"072C" => data_out<= x"B1";
        when x"072D" => data_out<= x"0C";
        when x"072E" => data_out<= x"C8";
        when x"072F" => data_out<= x"11";
        when x"0730" => data_out<= x"0C";
        when x"0731" => data_out<= x"D0";
        when x"0732" => data_out<= x"07";
        when x"0733" => data_out<= x"AA";
        when x"0734" => data_out<= x"A9";
        when x"0735" => data_out<= x"40";
        when x"0736" => data_out<= x"88";
        when x"0737" => data_out<= x"20";
        when x"0738" => data_out<= x"C5";
        when x"0739" => data_out<= x"B0";
        when x"073A" => data_out<= x"A0";
        when x"073B" => data_out<= x"14";
        when x"073C" => data_out<= x"20";
        when x"073D" => data_out<= x"93";
        when x"073E" => data_out<= x"B0";
        when x"073F" => data_out<= x"A0";
        when x"0740" => data_out<= x"12";
        when x"0741" => data_out<= x"20";
        when x"0742" => data_out<= x"4F";
        when x"0743" => data_out<= x"AF";
        when x"0744" => data_out<= x"20";
        when x"0745" => data_out<= x"6F";
        when x"0746" => data_out<= x"89";
        when x"0747" => data_out<= x"4C";
        when x"0748" => data_out<= x"41";
        when x"0749" => data_out<= x"89";
        when x"074A" => data_out<= x"C8";
        when x"074B" => data_out<= x"20";
        when x"074C" => data_out<= x"93";
        when x"074D" => data_out<= x"B0";
        when x"074E" => data_out<= x"A9";
        when x"074F" => data_out<= x"13";
        when x"0750" => data_out<= x"20";
        when x"0751" => data_out<= x"69";
        when x"0752" => data_out<= x"AF";
        when x"0753" => data_out<= x"20";
        when x"0754" => data_out<= x"50";
        when x"0755" => data_out<= x"8D";
        when x"0756" => data_out<= x"A0";
        when x"0757" => data_out<= x"13";
        when x"0758" => data_out<= x"20";
        when x"0759" => data_out<= x"C5";
        when x"075A" => data_out<= x"B0";
        when x"075B" => data_out<= x"A0";
        when x"075C" => data_out<= x"11";
        when x"075D" => data_out<= x"B1";
        when x"075E" => data_out<= x"0C";
        when x"075F" => data_out<= x"C8";
        when x"0760" => data_out<= x"11";
        when x"0761" => data_out<= x"0C";
        when x"0762" => data_out<= x"D0";
        when x"0763" => data_out<= x"0C";
        when x"0764" => data_out<= x"AD";
        when x"0765" => data_out<= x"00";
        when x"0766" => data_out<= x"02";
        when x"0767" => data_out<= x"AE";
        when x"0768" => data_out<= x"01";
        when x"0769" => data_out<= x"02";
        when x"076A" => data_out<= x"88";
        when x"076B" => data_out<= x"20";
        when x"076C" => data_out<= x"C5";
        when x"076D" => data_out<= x"B0";
        when x"076E" => data_out<= x"A0";
        when x"076F" => data_out<= x"12";
        when x"0770" => data_out<= x"20";
        when x"0771" => data_out<= x"4F";
        when x"0772" => data_out<= x"AF";
        when x"0773" => data_out<= x"20";
        when x"0774" => data_out<= x"D7";
        when x"0775" => data_out<= x"8D";
        when x"0776" => data_out<= x"4C";
        when x"0777" => data_out<= x"41";
        when x"0778" => data_out<= x"89";
        when x"0779" => data_out<= x"C8";
        when x"077A" => data_out<= x"20";
        when x"077B" => data_out<= x"93";
        when x"077C" => data_out<= x"B0";
        when x"077D" => data_out<= x"A9";
        when x"077E" => data_out<= x"13";
        when x"077F" => data_out<= x"20";
        when x"0780" => data_out<= x"69";
        when x"0781" => data_out<= x"AF";
        when x"0782" => data_out<= x"20";
        when x"0783" => data_out<= x"50";
        when x"0784" => data_out<= x"8D";
        when x"0785" => data_out<= x"A0";
        when x"0786" => data_out<= x"13";
        when x"0787" => data_out<= x"20";
        when x"0788" => data_out<= x"C5";
        when x"0789" => data_out<= x"B0";
        when x"078A" => data_out<= x"20";
        when x"078B" => data_out<= x"7B";
        when x"078C" => data_out<= x"B0";
        when x"078D" => data_out<= x"A9";
        when x"078E" => data_out<= x"11";
        when x"078F" => data_out<= x"20";
        when x"0790" => data_out<= x"69";
        when x"0791" => data_out<= x"AF";
        when x"0792" => data_out<= x"20";
        when x"0793" => data_out<= x"50";
        when x"0794" => data_out<= x"8D";
        when x"0795" => data_out<= x"A0";
        when x"0796" => data_out<= x"13";
        when x"0797" => data_out<= x"20";
        when x"0798" => data_out<= x"C5";
        when x"0799" => data_out<= x"B0";
        when x"079A" => data_out<= x"20";
        when x"079B" => data_out<= x"7B";
        when x"079C" => data_out<= x"B0";
        when x"079D" => data_out<= x"A9";
        when x"079E" => data_out<= x"0F";
        when x"079F" => data_out<= x"20";
        when x"07A0" => data_out<= x"69";
        when x"07A1" => data_out<= x"AF";
        when x"07A2" => data_out<= x"20";
        when x"07A3" => data_out<= x"50";
        when x"07A4" => data_out<= x"8D";
        when x"07A5" => data_out<= x"A0";
        when x"07A6" => data_out<= x"13";
        when x"07A7" => data_out<= x"20";
        when x"07A8" => data_out<= x"C5";
        when x"07A9" => data_out<= x"B0";
        when x"07AA" => data_out<= x"A0";
        when x"07AB" => data_out<= x"14";
        when x"07AC" => data_out<= x"20";
        when x"07AD" => data_out<= x"93";
        when x"07AE" => data_out<= x"B0";
        when x"07AF" => data_out<= x"A0";
        when x"07B0" => data_out<= x"14";
        when x"07B1" => data_out<= x"20";
        when x"07B2" => data_out<= x"93";
        when x"07B3" => data_out<= x"B0";
        when x"07B4" => data_out<= x"A0";
        when x"07B5" => data_out<= x"11";
        when x"07B6" => data_out<= x"B1";
        when x"07B7" => data_out<= x"0C";
        when x"07B8" => data_out<= x"20";
        when x"07B9" => data_out<= x"DF";
        when x"07BA" => data_out<= x"8A";
        when x"07BB" => data_out<= x"A9";
        when x"07BC" => data_out<= x"13";
        when x"07BD" => data_out<= x"A2";
        when x"07BE" => data_out<= x"BC";
        when x"07BF" => data_out<= x"20";
        when x"07C0" => data_out<= x"22";
        when x"07C1" => data_out<= x"81";
        when x"07C2" => data_out<= x"A0";
        when x"07C3" => data_out<= x"12";
        when x"07C4" => data_out<= x"20";
        when x"07C5" => data_out<= x"4F";
        when x"07C6" => data_out<= x"AF";
        when x"07C7" => data_out<= x"20";
        when x"07C8" => data_out<= x"31";
        when x"07C9" => data_out<= x"8C";
        when x"07CA" => data_out<= x"A9";
        when x"07CB" => data_out<= x"7D";
        when x"07CC" => data_out<= x"A2";
        when x"07CD" => data_out<= x"BD";
        when x"07CE" => data_out<= x"20";
        when x"07CF" => data_out<= x"22";
        when x"07D0" => data_out<= x"81";
        when x"07D1" => data_out<= x"A0";
        when x"07D2" => data_out<= x"10";
        when x"07D3" => data_out<= x"20";
        when x"07D4" => data_out<= x"4F";
        when x"07D5" => data_out<= x"AF";
        when x"07D6" => data_out<= x"18";
        when x"07D7" => data_out<= x"A0";
        when x"07D8" => data_out<= x"11";
        when x"07D9" => data_out<= x"71";
        when x"07DA" => data_out<= x"0C";
        when x"07DB" => data_out<= x"48";
        when x"07DC" => data_out<= x"8A";
        when x"07DD" => data_out<= x"C8";
        when x"07DE" => data_out<= x"71";
        when x"07DF" => data_out<= x"0C";
        when x"07E0" => data_out<= x"AA";
        when x"07E1" => data_out<= x"68";
        when x"07E2" => data_out<= x"20";
        when x"07E3" => data_out<= x"5A";
        when x"07E4" => data_out<= x"AE";
        when x"07E5" => data_out<= x"20";
        when x"07E6" => data_out<= x"31";
        when x"07E7" => data_out<= x"8C";
        when x"07E8" => data_out<= x"A9";
        when x"07E9" => data_out<= x"42";
        when x"07EA" => data_out<= x"A2";
        when x"07EB" => data_out<= x"BC";
        when x"07EC" => data_out<= x"20";
        when x"07ED" => data_out<= x"22";
        when x"07EE" => data_out<= x"81";
        when x"07EF" => data_out<= x"A0";
        when x"07F0" => data_out<= x"0D";
        when x"07F1" => data_out<= x"B1";
        when x"07F2" => data_out<= x"0C";
        when x"07F3" => data_out<= x"20";
        when x"07F4" => data_out<= x"FD";
        when x"07F5" => data_out<= x"8B";
        when x"07F6" => data_out<= x"20";
        when x"07F7" => data_out<= x"45";
        when x"07F8" => data_out<= x"8C";
        when x"07F9" => data_out<= x"4C";
        when x"07FA" => data_out<= x"41";
        when x"07FB" => data_out<= x"89";
        when x"07FC" => data_out<= x"C8";
        when x"07FD" => data_out<= x"20";
        when x"07FE" => data_out<= x"93";
        when x"07FF" => data_out<= x"B0";
        when x"0800" => data_out<= x"A9";
        when x"0801" => data_out<= x"13";
        when x"0802" => data_out<= x"20";
        when x"0803" => data_out<= x"69";
        when x"0804" => data_out<= x"AF";
        when x"0805" => data_out<= x"20";
        when x"0806" => data_out<= x"50";
        when x"0807" => data_out<= x"8D";
        when x"0808" => data_out<= x"A0";
        when x"0809" => data_out<= x"13";
        when x"080A" => data_out<= x"20";
        when x"080B" => data_out<= x"C5";
        when x"080C" => data_out<= x"B0";
        when x"080D" => data_out<= x"A0";
        when x"080E" => data_out<= x"11";
        when x"080F" => data_out<= x"B1";
        when x"0810" => data_out<= x"0C";
        when x"0811" => data_out<= x"C8";
        when x"0812" => data_out<= x"11";
        when x"0813" => data_out<= x"0C";
        when x"0814" => data_out<= x"D0";
        when x"0815" => data_out<= x"0A";
        when x"0816" => data_out<= x"AD";
        when x"0817" => data_out<= x"00";
        when x"0818" => data_out<= x"02";
        when x"0819" => data_out<= x"AE";
        when x"081A" => data_out<= x"01";
        when x"081B" => data_out<= x"02";
        when x"081C" => data_out<= x"88";
        when x"081D" => data_out<= x"20";
        when x"081E" => data_out<= x"C5";
        when x"081F" => data_out<= x"B0";
        when x"0820" => data_out<= x"A0";
        when x"0821" => data_out<= x"16";
        when x"0822" => data_out<= x"20";
        when x"0823" => data_out<= x"93";
        when x"0824" => data_out<= x"B0";
        when x"0825" => data_out<= x"A9";
        when x"0826" => data_out<= x"11";
        when x"0827" => data_out<= x"20";
        when x"0828" => data_out<= x"69";
        when x"0829" => data_out<= x"AF";
        when x"082A" => data_out<= x"20";
        when x"082B" => data_out<= x"50";
        when x"082C" => data_out<= x"8D";
        when x"082D" => data_out<= x"A0";
        when x"082E" => data_out<= x"13";
        when x"082F" => data_out<= x"20";
        when x"0830" => data_out<= x"C5";
        when x"0831" => data_out<= x"B0";
        when x"0832" => data_out<= x"A0";
        when x"0833" => data_out<= x"0F";
        when x"0834" => data_out<= x"B1";
        when x"0835" => data_out<= x"0C";
        when x"0836" => data_out<= x"C8";
        when x"0837" => data_out<= x"11";
        when x"0838" => data_out<= x"0C";
        when x"0839" => data_out<= x"D0";
        when x"083A" => data_out<= x"07";
        when x"083B" => data_out<= x"AA";
        when x"083C" => data_out<= x"98";
        when x"083D" => data_out<= x"88";
        when x"083E" => data_out<= x"20";
        when x"083F" => data_out<= x"C5";
        when x"0840" => data_out<= x"B0";
        when x"0841" => data_out<= x"A8";
        when x"0842" => data_out<= x"20";
        when x"0843" => data_out<= x"4F";
        when x"0844" => data_out<= x"AF";
        when x"0845" => data_out<= x"C9";
        when x"0846" => data_out<= x"00";
        when x"0847" => data_out<= x"8A";
        when x"0848" => data_out<= x"E9";
        when x"0849" => data_out<= x"01";
        when x"084A" => data_out<= x"90";
        when x"084B" => data_out<= x"13";
        when x"084C" => data_out<= x"A9";
        when x"084D" => data_out<= x"C0";
        when x"084E" => data_out<= x"A2";
        when x"084F" => data_out<= x"B9";
        when x"0850" => data_out<= x"20";
        when x"0851" => data_out<= x"22";
        when x"0852" => data_out<= x"81";
        when x"0853" => data_out<= x"20";
        when x"0854" => data_out<= x"45";
        when x"0855" => data_out<= x"8C";
        when x"0856" => data_out<= x"A2";
        when x"0857" => data_out<= x"00";
        when x"0858" => data_out<= x"A9";
        when x"0859" => data_out<= x"FF";
        when x"085A" => data_out<= x"A0";
        when x"085B" => data_out<= x"0F";
        when x"085C" => data_out<= x"20";
        when x"085D" => data_out<= x"C5";
        when x"085E" => data_out<= x"B0";
        when x"085F" => data_out<= x"A0";
        when x"0860" => data_out<= x"14";
        when x"0861" => data_out<= x"20";
        when x"0862" => data_out<= x"93";
        when x"0863" => data_out<= x"B0";
        when x"0864" => data_out<= x"A0";
        when x"0865" => data_out<= x"11";
        when x"0866" => data_out<= x"B1";
        when x"0867" => data_out<= x"0C";
        when x"0868" => data_out<= x"20";
        when x"0869" => data_out<= x"78";
        when x"086A" => data_out<= x"92";
        when x"086B" => data_out<= x"4C";
        when x"086C" => data_out<= x"41";
        when x"086D" => data_out<= x"89";
        when x"086E" => data_out<= x"20";
        when x"086F" => data_out<= x"1C";
        when x"0870" => data_out<= x"94";
        when x"0871" => data_out<= x"4C";
        when x"0872" => data_out<= x"41";
        when x"0873" => data_out<= x"89";
        when x"0874" => data_out<= x"A9";
        when x"0875" => data_out<= x"ED";
        when x"0876" => data_out<= x"A2";
        when x"0877" => data_out<= x"B4";
        when x"0878" => data_out<= x"20";
        when x"0879" => data_out<= x"22";
        when x"087A" => data_out<= x"81";
        when x"087B" => data_out<= x"4C";
        when x"087C" => data_out<= x"41";
        when x"087D" => data_out<= x"89";
        when x"087E" => data_out<= x"A9";
        when x"087F" => data_out<= x"3E";
        when x"0880" => data_out<= x"A2";
        when x"0881" => data_out<= x"B8";
        when x"0882" => data_out<= x"20";
        when x"0883" => data_out<= x"22";
        when x"0884" => data_out<= x"81";
        when x"0885" => data_out<= x"20";
        when x"0886" => data_out<= x"45";
        when x"0887" => data_out<= x"8C";
        when x"0888" => data_out<= x"A2";
        when x"0889" => data_out<= x"00";
        when x"088A" => data_out<= x"A9";
        when x"088B" => data_out<= x"02";
        when x"088C" => data_out<= x"4C";
        when x"088D" => data_out<= x"44";
        when x"088E" => data_out<= x"89";
        when x"088F" => data_out<= x"A0";
        when x"0890" => data_out<= x"14";
        when x"0891" => data_out<= x"20";
        when x"0892" => data_out<= x"4F";
        when x"0893" => data_out<= x"AF";
        when x"0894" => data_out<= x"20";
        when x"0895" => data_out<= x"E2";
        when x"0896" => data_out<= x"AE";
        when x"0897" => data_out<= x"A0";
        when x"0898" => data_out<= x"13";
        when x"0899" => data_out<= x"20";
        when x"089A" => data_out<= x"C5";
        when x"089B" => data_out<= x"B0";
        when x"089C" => data_out<= x"A0";
        when x"089D" => data_out<= x"14";
        when x"089E" => data_out<= x"20";
        when x"089F" => data_out<= x"4F";
        when x"08A0" => data_out<= x"AF";
        when x"08A1" => data_out<= x"85";
        when x"08A2" => data_out<= x"14";
        when x"08A3" => data_out<= x"86";
        when x"08A4" => data_out<= x"15";
        when x"08A5" => data_out<= x"A0";
        when x"08A6" => data_out<= x"00";
        when x"08A7" => data_out<= x"B1";
        when x"08A8" => data_out<= x"14";
        when x"08A9" => data_out<= x"C9";
        when x"08AA" => data_out<= x"20";
        when x"08AB" => data_out<= x"F0";
        when x"08AC" => data_out<= x"E2";
        when x"08AD" => data_out<= x"A0";
        when x"08AE" => data_out<= x"14";
        when x"08AF" => data_out<= x"20";
        when x"08B0" => data_out<= x"4F";
        when x"08B1" => data_out<= x"AF";
        when x"08B2" => data_out<= x"85";
        when x"08B3" => data_out<= x"14";
        when x"08B4" => data_out<= x"86";
        when x"08B5" => data_out<= x"15";
        when x"08B6" => data_out<= x"A0";
        when x"08B7" => data_out<= x"00";
        when x"08B8" => data_out<= x"B1";
        when x"08B9" => data_out<= x"14";
        when x"08BA" => data_out<= x"D0";
        when x"08BB" => data_out<= x"06";
        when x"08BC" => data_out<= x"20";
        when x"08BD" => data_out<= x"99";
        when x"08BE" => data_out<= x"9B";
        when x"08BF" => data_out<= x"4C";
        when x"08C0" => data_out<= x"41";
        when x"08C1" => data_out<= x"89";
        when x"08C2" => data_out<= x"A0";
        when x"08C3" => data_out<= x"16";
        when x"08C4" => data_out<= x"20";
        when x"08C5" => data_out<= x"93";
        when x"08C6" => data_out<= x"B0";
        when x"08C7" => data_out<= x"A9";
        when x"08C8" => data_out<= x"3F";
        when x"08C9" => data_out<= x"A2";
        when x"08CA" => data_out<= x"B6";
        when x"08CB" => data_out<= x"20";
        when x"08CC" => data_out<= x"F9";
        when x"08CD" => data_out<= x"9A";
        when x"08CE" => data_out<= x"AA";
        when x"08CF" => data_out<= x"D0";
        when x"08D0" => data_out<= x"4B";
        when x"08D1" => data_out<= x"A0";
        when x"08D2" => data_out<= x"16";
        when x"08D3" => data_out<= x"20";
        when x"08D4" => data_out<= x"93";
        when x"08D5" => data_out<= x"B0";
        when x"08D6" => data_out<= x"A9";
        when x"08D7" => data_out<= x"80";
        when x"08D8" => data_out<= x"A2";
        when x"08D9" => data_out<= x"BD";
        when x"08DA" => data_out<= x"20";
        when x"08DB" => data_out<= x"F9";
        when x"08DC" => data_out<= x"9A";
        when x"08DD" => data_out<= x"AA";
        when x"08DE" => data_out<= x"D0";
        when x"08DF" => data_out<= x"3C";
        when x"08E0" => data_out<= x"A0";
        when x"08E1" => data_out<= x"16";
        when x"08E2" => data_out<= x"20";
        when x"08E3" => data_out<= x"93";
        when x"08E4" => data_out<= x"B0";
        when x"08E5" => data_out<= x"A9";
        when x"08E6" => data_out<= x"9A";
        when x"08E7" => data_out<= x"A2";
        when x"08E8" => data_out<= x"BC";
        when x"08E9" => data_out<= x"20";
        when x"08EA" => data_out<= x"F9";
        when x"08EB" => data_out<= x"9A";
        when x"08EC" => data_out<= x"AA";
        when x"08ED" => data_out<= x"D0";
        when x"08EE" => data_out<= x"2D";
        when x"08EF" => data_out<= x"A0";
        when x"08F0" => data_out<= x"16";
        when x"08F1" => data_out<= x"20";
        when x"08F2" => data_out<= x"93";
        when x"08F3" => data_out<= x"B0";
        when x"08F4" => data_out<= x"A9";
        when x"08F5" => data_out<= x"95";
        when x"08F6" => data_out<= x"A2";
        when x"08F7" => data_out<= x"BC";
        when x"08F8" => data_out<= x"20";
        when x"08F9" => data_out<= x"F9";
        when x"08FA" => data_out<= x"9A";
        when x"08FB" => data_out<= x"AA";
        when x"08FC" => data_out<= x"D0";
        when x"08FD" => data_out<= x"1E";
        when x"08FE" => data_out<= x"A0";
        when x"08FF" => data_out<= x"16";
        when x"0900" => data_out<= x"20";
        when x"0901" => data_out<= x"93";
        when x"0902" => data_out<= x"B0";
        when x"0903" => data_out<= x"A9";
        when x"0904" => data_out<= x"11";
        when x"0905" => data_out<= x"A2";
        when x"0906" => data_out<= x"BD";
        when x"0907" => data_out<= x"20";
        when x"0908" => data_out<= x"F9";
        when x"0909" => data_out<= x"9A";
        when x"090A" => data_out<= x"AA";
        when x"090B" => data_out<= x"D0";
        when x"090C" => data_out<= x"0F";
        when x"090D" => data_out<= x"A0";
        when x"090E" => data_out<= x"16";
        when x"090F" => data_out<= x"20";
        when x"0910" => data_out<= x"93";
        when x"0911" => data_out<= x"B0";
        when x"0912" => data_out<= x"A9";
        when x"0913" => data_out<= x"39";
        when x"0914" => data_out<= x"A2";
        when x"0915" => data_out<= x"BD";
        when x"0916" => data_out<= x"20";
        when x"0917" => data_out<= x"F9";
        when x"0918" => data_out<= x"9A";
        when x"0919" => data_out<= x"AA";
        when x"091A" => data_out<= x"F0";
        when x"091B" => data_out<= x"0B";
        when x"091C" => data_out<= x"A0";
        when x"091D" => data_out<= x"14";
        when x"091E" => data_out<= x"20";
        when x"091F" => data_out<= x"4F";
        when x"0920" => data_out<= x"AF";
        when x"0921" => data_out<= x"20";
        when x"0922" => data_out<= x"F4";
        when x"0923" => data_out<= x"9C";
        when x"0924" => data_out<= x"4C";
        when x"0925" => data_out<= x"41";
        when x"0926" => data_out<= x"89";
        when x"0927" => data_out<= x"A0";
        when x"0928" => data_out<= x"14";
        when x"0929" => data_out<= x"20";
        when x"092A" => data_out<= x"4F";
        when x"092B" => data_out<= x"AF";
        when x"092C" => data_out<= x"85";
        when x"092D" => data_out<= x"14";
        when x"092E" => data_out<= x"86";
        when x"092F" => data_out<= x"15";
        when x"0930" => data_out<= x"A0";
        when x"0931" => data_out<= x"00";
        when x"0932" => data_out<= x"B1";
        when x"0933" => data_out<= x"14";
        when x"0934" => data_out<= x"20";
        when x"0935" => data_out<= x"05";
        when x"0936" => data_out<= x"9C";
        when x"0937" => data_out<= x"4C";
        when x"0938" => data_out<= x"41";
        when x"0939" => data_out<= x"89";
        when x"093A" => data_out<= x"A9";
        when x"093B" => data_out<= x"62";
        when x"093C" => data_out<= x"A2";
        when x"093D" => data_out<= x"B5";
        when x"093E" => data_out<= x"20";
        when x"093F" => data_out<= x"99";
        when x"0940" => data_out<= x"8C";
        when x"0941" => data_out<= x"A2";
        when x"0942" => data_out<= x"00";
        when x"0943" => data_out<= x"8A";
        when x"0944" => data_out<= x"A0";
        when x"0945" => data_out<= x"18";
        when x"0946" => data_out<= x"4C";
        when x"0947" => data_out<= x"14";
        when x"0948" => data_out<= x"AE";
        when x"0949" => data_out<= x"20";
        when x"094A" => data_out<= x"7B";
        when x"094B" => data_out<= x"B0";
        when x"094C" => data_out<= x"20";
        when x"094D" => data_out<= x"4D";
        when x"094E" => data_out<= x"AF";
        when x"094F" => data_out<= x"85";
        when x"0950" => data_out<= x"14";
        when x"0951" => data_out<= x"86";
        when x"0952" => data_out<= x"15";
        when x"0953" => data_out<= x"A2";
        when x"0954" => data_out<= x"00";
        when x"0955" => data_out<= x"A1";
        when x"0956" => data_out<= x"14";
        when x"0957" => data_out<= x"4C";
        when x"0958" => data_out<= x"14";
        when x"0959" => data_out<= x"AF";
        when x"095A" => data_out<= x"20";
        when x"095B" => data_out<= x"65";
        when x"095C" => data_out<= x"B0";
        when x"095D" => data_out<= x"A0";
        when x"095E" => data_out<= x"02";
        when x"095F" => data_out<= x"20";
        when x"0960" => data_out<= x"4F";
        when x"0961" => data_out<= x"AF";
        when x"0962" => data_out<= x"85";
        when x"0963" => data_out<= x"14";
        when x"0964" => data_out<= x"86";
        when x"0965" => data_out<= x"15";
        when x"0966" => data_out<= x"A0";
        when x"0967" => data_out<= x"00";
        when x"0968" => data_out<= x"B1";
        when x"0969" => data_out<= x"0C";
        when x"096A" => data_out<= x"91";
        when x"096B" => data_out<= x"14";
        when x"096C" => data_out<= x"4C";
        when x"096D" => data_out<= x"22";
        when x"096E" => data_out<= x"AF";
        when x"096F" => data_out<= x"20";
        when x"0970" => data_out<= x"7B";
        when x"0971" => data_out<= x"B0";
        when x"0972" => data_out<= x"A0";
        when x"0973" => data_out<= x"15";
        when x"0974" => data_out<= x"20";
        when x"0975" => data_out<= x"13";
        when x"0976" => data_out<= x"B1";
        when x"0977" => data_out<= x"A2";
        when x"0978" => data_out<= x"00";
        when x"0979" => data_out<= x"8A";
        when x"097A" => data_out<= x"A0";
        when x"097B" => data_out<= x"13";
        when x"097C" => data_out<= x"20";
        when x"097D" => data_out<= x"C5";
        when x"097E" => data_out<= x"B0";
        when x"097F" => data_out<= x"A0";
        when x"0980" => data_out<= x"14";
        when x"0981" => data_out<= x"20";
        when x"0982" => data_out<= x"4F";
        when x"0983" => data_out<= x"AF";
        when x"0984" => data_out<= x"A0";
        when x"0985" => data_out<= x"15";
        when x"0986" => data_out<= x"D1";
        when x"0987" => data_out<= x"0C";
        when x"0988" => data_out<= x"8A";
        when x"0989" => data_out<= x"C8";
        when x"098A" => data_out<= x"F1";
        when x"098B" => data_out<= x"0C";
        when x"098C" => data_out<= x"90";
        when x"098D" => data_out<= x"03";
        when x"098E" => data_out<= x"4C";
        when x"098F" => data_out<= x"C9";
        when x"0990" => data_out<= x"8A";
        when x"0991" => data_out<= x"A0";
        when x"0992" => data_out<= x"14";
        when x"0993" => data_out<= x"20";
        when x"0994" => data_out<= x"4F";
        when x"0995" => data_out<= x"AF";
        when x"0996" => data_out<= x"18";
        when x"0997" => data_out<= x"A0";
        when x"0998" => data_out<= x"17";
        when x"0999" => data_out<= x"71";
        when x"099A" => data_out<= x"0C";
        when x"099B" => data_out<= x"48";
        when x"099C" => data_out<= x"8A";
        when x"099D" => data_out<= x"C8";
        when x"099E" => data_out<= x"71";
        when x"099F" => data_out<= x"0C";
        when x"09A0" => data_out<= x"AA";
        when x"09A1" => data_out<= x"68";
        when x"09A2" => data_out<= x"20";
        when x"09A3" => data_out<= x"C3";
        when x"09A4" => data_out<= x"B0";
        when x"09A5" => data_out<= x"20";
        when x"09A6" => data_out<= x"31";
        when x"09A7" => data_out<= x"8C";
        when x"09A8" => data_out<= x"A9";
        when x"09A9" => data_out<= x"99";
        when x"09AA" => data_out<= x"A2";
        when x"09AB" => data_out<= x"B5";
        when x"09AC" => data_out<= x"20";
        when x"09AD" => data_out<= x"22";
        when x"09AE" => data_out<= x"81";
        when x"09AF" => data_out<= x"A9";
        when x"09B0" => data_out<= x"00";
        when x"09B1" => data_out<= x"A0";
        when x"09B2" => data_out<= x"12";
        when x"09B3" => data_out<= x"91";
        when x"09B4" => data_out<= x"0C";
        when x"09B5" => data_out<= x"C9";
        when x"09B6" => data_out<= x"10";
        when x"09B7" => data_out<= x"B0";
        when x"09B8" => data_out<= x"77";
        when x"09B9" => data_out<= x"B1";
        when x"09BA" => data_out<= x"0C";
        when x"09BB" => data_out<= x"18";
        when x"09BC" => data_out<= x"C8";
        when x"09BD" => data_out<= x"71";
        when x"09BE" => data_out<= x"0C";
        when x"09BF" => data_out<= x"48";
        when x"09C0" => data_out<= x"A9";
        when x"09C1" => data_out<= x"00";
        when x"09C2" => data_out<= x"C8";
        when x"09C3" => data_out<= x"71";
        when x"09C4" => data_out<= x"0C";
        when x"09C5" => data_out<= x"AA";
        when x"09C6" => data_out<= x"68";
        when x"09C7" => data_out<= x"C8";
        when x"09C8" => data_out<= x"D1";
        when x"09C9" => data_out<= x"0C";
        when x"09CA" => data_out<= x"8A";
        when x"09CB" => data_out<= x"C8";
        when x"09CC" => data_out<= x"F1";
        when x"09CD" => data_out<= x"0C";
        when x"09CE" => data_out<= x"B0";
        when x"09CF" => data_out<= x"5E";
        when x"09D0" => data_out<= x"A9";
        when x"09D1" => data_out<= x"02";
        when x"09D2" => data_out<= x"20";
        when x"09D3" => data_out<= x"69";
        when x"09D4" => data_out<= x"AF";
        when x"09D5" => data_out<= x"A0";
        when x"09D6" => data_out<= x"12";
        when x"09D7" => data_out<= x"18";
        when x"09D8" => data_out<= x"71";
        when x"09D9" => data_out<= x"0C";
        when x"09DA" => data_out<= x"90";
        when x"09DB" => data_out<= x"01";
        when x"09DC" => data_out<= x"E8";
        when x"09DD" => data_out<= x"20";
        when x"09DE" => data_out<= x"7B";
        when x"09DF" => data_out<= x"B0";
        when x"09E0" => data_out<= x"A0";
        when x"09E1" => data_out<= x"14";
        when x"09E2" => data_out<= x"B1";
        when x"09E3" => data_out<= x"0C";
        when x"09E4" => data_out<= x"18";
        when x"09E5" => data_out<= x"A0";
        when x"09E6" => data_out<= x"02";
        when x"09E7" => data_out<= x"71";
        when x"09E8" => data_out<= x"0C";
        when x"09E9" => data_out<= x"48";
        when x"09EA" => data_out<= x"A9";
        when x"09EB" => data_out<= x"00";
        when x"09EC" => data_out<= x"C8";
        when x"09ED" => data_out<= x"71";
        when x"09EE" => data_out<= x"0C";
        when x"09EF" => data_out<= x"AA";
        when x"09F0" => data_out<= x"68";
        when x"09F1" => data_out<= x"20";
        when x"09F2" => data_out<= x"49";
        when x"09F3" => data_out<= x"89";
        when x"09F4" => data_out<= x"A0";
        when x"09F5" => data_out<= x"00";
        when x"09F6" => data_out<= x"20";
        when x"09F7" => data_out<= x"AD";
        when x"09F8" => data_out<= x"B0";
        when x"09F9" => data_out<= x"A9";
        when x"09FA" => data_out<= x"02";
        when x"09FB" => data_out<= x"20";
        when x"09FC" => data_out<= x"69";
        when x"09FD" => data_out<= x"AF";
        when x"09FE" => data_out<= x"A0";
        when x"09FF" => data_out<= x"12";
        when x"0A00" => data_out<= x"18";
        when x"0A01" => data_out<= x"71";
        when x"0A02" => data_out<= x"0C";
        when x"0A03" => data_out<= x"90";
        when x"0A04" => data_out<= x"01";
        when x"0A05" => data_out<= x"E8";
        when x"0A06" => data_out<= x"85";
        when x"0A07" => data_out<= x"14";
        when x"0A08" => data_out<= x"86";
        when x"0A09" => data_out<= x"15";
        when x"0A0A" => data_out<= x"A0";
        when x"0A0B" => data_out<= x"00";
        when x"0A0C" => data_out<= x"B1";
        when x"0A0D" => data_out<= x"14";
        when x"0A0E" => data_out<= x"20";
        when x"0A0F" => data_out<= x"FD";
        when x"0A10" => data_out<= x"8B";
        when x"0A11" => data_out<= x"20";
        when x"0A12" => data_out<= x"8C";
        when x"0A13" => data_out<= x"8C";
        when x"0A14" => data_out<= x"A0";
        when x"0A15" => data_out<= x"12";
        when x"0A16" => data_out<= x"B1";
        when x"0A17" => data_out<= x"0C";
        when x"0A18" => data_out<= x"18";
        when x"0A19" => data_out<= x"69";
        when x"0A1A" => data_out<= x"01";
        when x"0A1B" => data_out<= x"4C";
        when x"0A1C" => data_out<= x"B3";
        when x"0A1D" => data_out<= x"89";
        when x"0A1E" => data_out<= x"A9";
        when x"0A1F" => data_out<= x"01";
        when x"0A20" => data_out<= x"A2";
        when x"0A21" => data_out<= x"BD";
        when x"0A22" => data_out<= x"20";
        when x"0A23" => data_out<= x"22";
        when x"0A24" => data_out<= x"81";
        when x"0A25" => data_out<= x"A0";
        when x"0A26" => data_out<= x"12";
        when x"0A27" => data_out<= x"B1";
        when x"0A28" => data_out<= x"0C";
        when x"0A29" => data_out<= x"18";
        when x"0A2A" => data_out<= x"69";
        when x"0A2B" => data_out<= x"01";
        when x"0A2C" => data_out<= x"91";
        when x"0A2D" => data_out<= x"0C";
        when x"0A2E" => data_out<= x"A0";
        when x"0A2F" => data_out<= x"12";
        when x"0A30" => data_out<= x"B1";
        when x"0A31" => data_out<= x"0C";
        when x"0A32" => data_out<= x"C9";
        when x"0A33" => data_out<= x"10";
        when x"0A34" => data_out<= x"90";
        when x"0A35" => data_out<= x"E8";
        when x"0A36" => data_out<= x"A9";
        when x"0A37" => data_out<= x"7C";
        when x"0A38" => data_out<= x"20";
        when x"0A39" => data_out<= x"F0";
        when x"0A3A" => data_out<= x"80";
        when x"0A3B" => data_out<= x"A9";
        when x"0A3C" => data_out<= x"00";
        when x"0A3D" => data_out<= x"A0";
        when x"0A3E" => data_out<= x"12";
        when x"0A3F" => data_out<= x"91";
        when x"0A40" => data_out<= x"0C";
        when x"0A41" => data_out<= x"C9";
        when x"0A42" => data_out<= x"10";
        when x"0A43" => data_out<= x"B0";
        when x"0A44" => data_out<= x"70";
        when x"0A45" => data_out<= x"B1";
        when x"0A46" => data_out<= x"0C";
        when x"0A47" => data_out<= x"18";
        when x"0A48" => data_out<= x"C8";
        when x"0A49" => data_out<= x"71";
        when x"0A4A" => data_out<= x"0C";
        when x"0A4B" => data_out<= x"48";
        when x"0A4C" => data_out<= x"A9";
        when x"0A4D" => data_out<= x"00";
        when x"0A4E" => data_out<= x"C8";
        when x"0A4F" => data_out<= x"71";
        when x"0A50" => data_out<= x"0C";
        when x"0A51" => data_out<= x"AA";
        when x"0A52" => data_out<= x"68";
        when x"0A53" => data_out<= x"C8";
        when x"0A54" => data_out<= x"D1";
        when x"0A55" => data_out<= x"0C";
        when x"0A56" => data_out<= x"8A";
        when x"0A57" => data_out<= x"C8";
        when x"0A58" => data_out<= x"F1";
        when x"0A59" => data_out<= x"0C";
        when x"0A5A" => data_out<= x"B0";
        when x"0A5B" => data_out<= x"59";
        when x"0A5C" => data_out<= x"A9";
        when x"0A5D" => data_out<= x"02";
        when x"0A5E" => data_out<= x"20";
        when x"0A5F" => data_out<= x"69";
        when x"0A60" => data_out<= x"AF";
        when x"0A61" => data_out<= x"A0";
        when x"0A62" => data_out<= x"12";
        when x"0A63" => data_out<= x"18";
        when x"0A64" => data_out<= x"71";
        when x"0A65" => data_out<= x"0C";
        when x"0A66" => data_out<= x"90";
        when x"0A67" => data_out<= x"01";
        when x"0A68" => data_out<= x"E8";
        when x"0A69" => data_out<= x"85";
        when x"0A6A" => data_out<= x"14";
        when x"0A6B" => data_out<= x"86";
        when x"0A6C" => data_out<= x"15";
        when x"0A6D" => data_out<= x"A0";
        when x"0A6E" => data_out<= x"00";
        when x"0A6F" => data_out<= x"B1";
        when x"0A70" => data_out<= x"14";
        when x"0A71" => data_out<= x"C9";
        when x"0A72" => data_out<= x"20";
        when x"0A73" => data_out<= x"90";
        when x"0A74" => data_out<= x"31";
        when x"0A75" => data_out<= x"A9";
        when x"0A76" => data_out<= x"02";
        when x"0A77" => data_out<= x"20";
        when x"0A78" => data_out<= x"69";
        when x"0A79" => data_out<= x"AF";
        when x"0A7A" => data_out<= x"A0";
        when x"0A7B" => data_out<= x"12";
        when x"0A7C" => data_out<= x"18";
        when x"0A7D" => data_out<= x"71";
        when x"0A7E" => data_out<= x"0C";
        when x"0A7F" => data_out<= x"90";
        when x"0A80" => data_out<= x"01";
        when x"0A81" => data_out<= x"E8";
        when x"0A82" => data_out<= x"85";
        when x"0A83" => data_out<= x"14";
        when x"0A84" => data_out<= x"86";
        when x"0A85" => data_out<= x"15";
        when x"0A86" => data_out<= x"A0";
        when x"0A87" => data_out<= x"00";
        when x"0A88" => data_out<= x"B1";
        when x"0A89" => data_out<= x"14";
        when x"0A8A" => data_out<= x"C9";
        when x"0A8B" => data_out<= x"7F";
        when x"0A8C" => data_out<= x"B0";
        when x"0A8D" => data_out<= x"18";
        when x"0A8E" => data_out<= x"A9";
        when x"0A8F" => data_out<= x"02";
        when x"0A90" => data_out<= x"20";
        when x"0A91" => data_out<= x"69";
        when x"0A92" => data_out<= x"AF";
        when x"0A93" => data_out<= x"A0";
        when x"0A94" => data_out<= x"12";
        when x"0A95" => data_out<= x"18";
        when x"0A96" => data_out<= x"71";
        when x"0A97" => data_out<= x"0C";
        when x"0A98" => data_out<= x"90";
        when x"0A99" => data_out<= x"01";
        when x"0A9A" => data_out<= x"E8";
        when x"0A9B" => data_out<= x"85";
        when x"0A9C" => data_out<= x"14";
        when x"0A9D" => data_out<= x"86";
        when x"0A9E" => data_out<= x"15";
        when x"0A9F" => data_out<= x"A0";
        when x"0AA0" => data_out<= x"00";
        when x"0AA1" => data_out<= x"B1";
        when x"0AA2" => data_out<= x"14";
        when x"0AA3" => data_out<= x"4C";
        when x"0AA4" => data_out<= x"A8";
        when x"0AA5" => data_out<= x"8A";
        when x"0AA6" => data_out<= x"A9";
        when x"0AA7" => data_out<= x"2E";
        when x"0AA8" => data_out<= x"20";
        when x"0AA9" => data_out<= x"F0";
        when x"0AAA" => data_out<= x"80";
        when x"0AAB" => data_out<= x"A0";
        when x"0AAC" => data_out<= x"12";
        when x"0AAD" => data_out<= x"B1";
        when x"0AAE" => data_out<= x"0C";
        when x"0AAF" => data_out<= x"18";
        when x"0AB0" => data_out<= x"69";
        when x"0AB1" => data_out<= x"01";
        when x"0AB2" => data_out<= x"4C";
        when x"0AB3" => data_out<= x"3F";
        when x"0AB4" => data_out<= x"8A";
        when x"0AB5" => data_out<= x"A9";
        when x"0AB6" => data_out<= x"7C";
        when x"0AB7" => data_out<= x"20";
        when x"0AB8" => data_out<= x"F0";
        when x"0AB9" => data_out<= x"80";
        when x"0ABA" => data_out<= x"20";
        when x"0ABB" => data_out<= x"45";
        when x"0ABC" => data_out<= x"8C";
        when x"0ABD" => data_out<= x"A0";
        when x"0ABE" => data_out<= x"13";
        when x"0ABF" => data_out<= x"A2";
        when x"0AC0" => data_out<= x"00";
        when x"0AC1" => data_out<= x"A9";
        when x"0AC2" => data_out<= x"10";
        when x"0AC3" => data_out<= x"20";
        when x"0AC4" => data_out<= x"04";
        when x"0AC5" => data_out<= x"AE";
        when x"0AC6" => data_out<= x"4C";
        when x"0AC7" => data_out<= x"7F";
        when x"0AC8" => data_out<= x"89";
        when x"0AC9" => data_out<= x"20";
        when x"0ACA" => data_out<= x"4F";
        when x"0ACB" => data_out<= x"AF";
        when x"0ACC" => data_out<= x"18";
        when x"0ACD" => data_out<= x"A0";
        when x"0ACE" => data_out<= x"17";
        when x"0ACF" => data_out<= x"71";
        when x"0AD0" => data_out<= x"0C";
        when x"0AD1" => data_out<= x"8D";
        when x"0AD2" => data_out<= x"00";
        when x"0AD3" => data_out<= x"02";
        when x"0AD4" => data_out<= x"8A";
        when x"0AD5" => data_out<= x"C8";
        when x"0AD6" => data_out<= x"71";
        when x"0AD7" => data_out<= x"0C";
        when x"0AD8" => data_out<= x"8D";
        when x"0AD9" => data_out<= x"01";
        when x"0ADA" => data_out<= x"02";
        when x"0ADB" => data_out<= x"C8";
        when x"0ADC" => data_out<= x"4C";
        when x"0ADD" => data_out<= x"14";
        when x"0ADE" => data_out<= x"AE";
        when x"0ADF" => data_out<= x"20";
        when x"0AE0" => data_out<= x"65";
        when x"0AE1" => data_out<= x"B0";
        when x"0AE2" => data_out<= x"20";
        when x"0AE3" => data_out<= x"73";
        when x"0AE4" => data_out<= x"AE";
        when x"0AE5" => data_out<= x"A2";
        when x"0AE6" => data_out<= x"00";
        when x"0AE7" => data_out<= x"8A";
        when x"0AE8" => data_out<= x"20";
        when x"0AE9" => data_out<= x"C3";
        when x"0AEA" => data_out<= x"B0";
        when x"0AEB" => data_out<= x"A0";
        when x"0AEC" => data_out<= x"03";
        when x"0AED" => data_out<= x"D1";
        when x"0AEE" => data_out<= x"0C";
        when x"0AEF" => data_out<= x"8A";
        when x"0AF0" => data_out<= x"C8";
        when x"0AF1" => data_out<= x"F1";
        when x"0AF2" => data_out<= x"0C";
        when x"0AF3" => data_out<= x"B0";
        when x"0AF4" => data_out<= x"22";
        when x"0AF5" => data_out<= x"20";
        when x"0AF6" => data_out<= x"4D";
        when x"0AF7" => data_out<= x"AF";
        when x"0AF8" => data_out<= x"18";
        when x"0AF9" => data_out<= x"A0";
        when x"0AFA" => data_out<= x"05";
        when x"0AFB" => data_out<= x"71";
        when x"0AFC" => data_out<= x"0C";
        when x"0AFD" => data_out<= x"48";
        when x"0AFE" => data_out<= x"8A";
        when x"0AFF" => data_out<= x"C8";
        when x"0B00" => data_out<= x"71";
        when x"0B01" => data_out<= x"0C";
        when x"0B02" => data_out<= x"AA";
        when x"0B03" => data_out<= x"68";
        when x"0B04" => data_out<= x"20";
        when x"0B05" => data_out<= x"7B";
        when x"0B06" => data_out<= x"B0";
        when x"0B07" => data_out<= x"A0";
        when x"0B08" => data_out<= x"04";
        when x"0B09" => data_out<= x"B1";
        when x"0B0A" => data_out<= x"0C";
        when x"0B0B" => data_out<= x"20";
        when x"0B0C" => data_out<= x"5A";
        when x"0B0D" => data_out<= x"89";
        when x"0B0E" => data_out<= x"20";
        when x"0B0F" => data_out<= x"4D";
        when x"0B10" => data_out<= x"AF";
        when x"0B11" => data_out<= x"20";
        when x"0B12" => data_out<= x"E2";
        when x"0B13" => data_out<= x"AE";
        when x"0B14" => data_out<= x"4C";
        when x"0B15" => data_out<= x"E8";
        when x"0B16" => data_out<= x"8A";
        when x"0B17" => data_out<= x"4C";
        when x"0B18" => data_out<= x"36";
        when x"0B19" => data_out<= x"AF";
        when x"0B1A" => data_out<= x"20";
        when x"0B1B" => data_out<= x"7B";
        when x"0B1C" => data_out<= x"B0";
        when x"0B1D" => data_out<= x"20";
        when x"0B1E" => data_out<= x"77";
        when x"0B1F" => data_out<= x"B0";
        when x"0B20" => data_out<= x"20";
        when x"0B21" => data_out<= x"6A";
        when x"0B22" => data_out<= x"AE";
        when x"0B23" => data_out<= x"A0";
        when x"0B24" => data_out<= x"00";
        when x"0B25" => data_out<= x"91";
        when x"0B26" => data_out<= x"0C";
        when x"0B27" => data_out<= x"C9";
        when x"0B28" => data_out<= x"04";
        when x"0B29" => data_out<= x"B0";
        when x"0B2A" => data_out<= x"58";
        when x"0B2B" => data_out<= x"A0";
        when x"0B2C" => data_out<= x"04";
        when x"0B2D" => data_out<= x"20";
        when x"0B2E" => data_out<= x"4F";
        when x"0B2F" => data_out<= x"AF";
        when x"0B30" => data_out<= x"85";
        when x"0B31" => data_out<= x"14";
        when x"0B32" => data_out<= x"86";
        when x"0B33" => data_out<= x"15";
        when x"0B34" => data_out<= x"A0";
        when x"0B35" => data_out<= x"00";
        when x"0B36" => data_out<= x"B1";
        when x"0B37" => data_out<= x"0C";
        when x"0B38" => data_out<= x"A8";
        when x"0B39" => data_out<= x"B1";
        when x"0B3A" => data_out<= x"14";
        when x"0B3B" => data_out<= x"F0";
        when x"0B3C" => data_out<= x"46";
        when x"0B3D" => data_out<= x"A0";
        when x"0B3E" => data_out<= x"04";
        when x"0B3F" => data_out<= x"20";
        when x"0B40" => data_out<= x"4F";
        when x"0B41" => data_out<= x"AF";
        when x"0B42" => data_out<= x"85";
        when x"0B43" => data_out<= x"14";
        when x"0B44" => data_out<= x"86";
        when x"0B45" => data_out<= x"15";
        when x"0B46" => data_out<= x"A0";
        when x"0B47" => data_out<= x"00";
        when x"0B48" => data_out<= x"B1";
        when x"0B49" => data_out<= x"0C";
        when x"0B4A" => data_out<= x"A8";
        when x"0B4B" => data_out<= x"B1";
        when x"0B4C" => data_out<= x"14";
        when x"0B4D" => data_out<= x"20";
        when x"0B4E" => data_out<= x"0B";
        when x"0B4F" => data_out<= x"8D";
        when x"0B50" => data_out<= x"AA";
        when x"0B51" => data_out<= x"F0";
        when x"0B52" => data_out<= x"30";
        when x"0B53" => data_out<= x"A0";
        when x"0B54" => data_out<= x"02";
        when x"0B55" => data_out<= x"20";
        when x"0B56" => data_out<= x"4F";
        when x"0B57" => data_out<= x"AF";
        when x"0B58" => data_out<= x"20";
        when x"0B59" => data_out<= x"29";
        when x"0B5A" => data_out<= x"AE";
        when x"0B5B" => data_out<= x"20";
        when x"0B5C" => data_out<= x"7B";
        when x"0B5D" => data_out<= x"B0";
        when x"0B5E" => data_out<= x"A0";
        when x"0B5F" => data_out<= x"06";
        when x"0B60" => data_out<= x"20";
        when x"0B61" => data_out<= x"4F";
        when x"0B62" => data_out<= x"AF";
        when x"0B63" => data_out<= x"85";
        when x"0B64" => data_out<= x"14";
        when x"0B65" => data_out<= x"86";
        when x"0B66" => data_out<= x"15";
        when x"0B67" => data_out<= x"A0";
        when x"0B68" => data_out<= x"02";
        when x"0B69" => data_out<= x"B1";
        when x"0B6A" => data_out<= x"0C";
        when x"0B6B" => data_out<= x"A8";
        when x"0B6C" => data_out<= x"B1";
        when x"0B6D" => data_out<= x"14";
        when x"0B6E" => data_out<= x"20";
        when x"0B6F" => data_out<= x"AF";
        when x"0B70" => data_out<= x"8C";
        when x"0B71" => data_out<= x"20";
        when x"0B72" => data_out<= x"43";
        when x"0B73" => data_out<= x"B0";
        when x"0B74" => data_out<= x"A0";
        when x"0B75" => data_out<= x"01";
        when x"0B76" => data_out<= x"20";
        when x"0B77" => data_out<= x"C5";
        when x"0B78" => data_out<= x"B0";
        when x"0B79" => data_out<= x"A0";
        when x"0B7A" => data_out<= x"00";
        when x"0B7B" => data_out<= x"B1";
        when x"0B7C" => data_out<= x"0C";
        when x"0B7D" => data_out<= x"18";
        when x"0B7E" => data_out<= x"69";
        when x"0B7F" => data_out<= x"01";
        when x"0B80" => data_out<= x"4C";
        when x"0B81" => data_out<= x"25";
        when x"0B82" => data_out<= x"8B";
        when x"0B83" => data_out<= x"A0";
        when x"0B84" => data_out<= x"02";
        when x"0B85" => data_out<= x"20";
        when x"0B86" => data_out<= x"4F";
        when x"0B87" => data_out<= x"AF";
        when x"0B88" => data_out<= x"4C";
        when x"0B89" => data_out<= x"2C";
        when x"0B8A" => data_out<= x"AF";
        when x"0B8B" => data_out<= x"20";
        when x"0B8C" => data_out<= x"7B";
        when x"0B8D" => data_out<= x"B0";
        when x"0B8E" => data_out<= x"A9";
        when x"0B8F" => data_out<= x"00";
        when x"0B90" => data_out<= x"20";
        when x"0B91" => data_out<= x"65";
        when x"0B92" => data_out<= x"B0";
        when x"0B93" => data_out<= x"20";
        when x"0B94" => data_out<= x"6A";
        when x"0B95" => data_out<= x"AE";
        when x"0B96" => data_out<= x"A8";
        when x"0B97" => data_out<= x"91";
        when x"0B98" => data_out<= x"0C";
        when x"0B99" => data_out<= x"C9";
        when x"0B9A" => data_out<= x"02";
        when x"0B9B" => data_out<= x"B0";
        when x"0B9C" => data_out<= x"57";
        when x"0B9D" => data_out<= x"A0";
        when x"0B9E" => data_out<= x"03";
        when x"0B9F" => data_out<= x"20";
        when x"0BA0" => data_out<= x"4F";
        when x"0BA1" => data_out<= x"AF";
        when x"0BA2" => data_out<= x"85";
        when x"0BA3" => data_out<= x"14";
        when x"0BA4" => data_out<= x"86";
        when x"0BA5" => data_out<= x"15";
        when x"0BA6" => data_out<= x"A0";
        when x"0BA7" => data_out<= x"00";
        when x"0BA8" => data_out<= x"B1";
        when x"0BA9" => data_out<= x"0C";
        when x"0BAA" => data_out<= x"A8";
        when x"0BAB" => data_out<= x"B1";
        when x"0BAC" => data_out<= x"14";
        when x"0BAD" => data_out<= x"F0";
        when x"0BAE" => data_out<= x"45";
        when x"0BAF" => data_out<= x"A0";
        when x"0BB0" => data_out<= x"03";
        when x"0BB1" => data_out<= x"20";
        when x"0BB2" => data_out<= x"4F";
        when x"0BB3" => data_out<= x"AF";
        when x"0BB4" => data_out<= x"85";
        when x"0BB5" => data_out<= x"14";
        when x"0BB6" => data_out<= x"86";
        when x"0BB7" => data_out<= x"15";
        when x"0BB8" => data_out<= x"A0";
        when x"0BB9" => data_out<= x"00";
        when x"0BBA" => data_out<= x"B1";
        when x"0BBB" => data_out<= x"0C";
        when x"0BBC" => data_out<= x"A8";
        when x"0BBD" => data_out<= x"B1";
        when x"0BBE" => data_out<= x"14";
        when x"0BBF" => data_out<= x"20";
        when x"0BC0" => data_out<= x"0B";
        when x"0BC1" => data_out<= x"8D";
        when x"0BC2" => data_out<= x"AA";
        when x"0BC3" => data_out<= x"F0";
        when x"0BC4" => data_out<= x"2F";
        when x"0BC5" => data_out<= x"A0";
        when x"0BC6" => data_out<= x"01";
        when x"0BC7" => data_out<= x"A2";
        when x"0BC8" => data_out<= x"00";
        when x"0BC9" => data_out<= x"B1";
        when x"0BCA" => data_out<= x"0C";
        when x"0BCB" => data_out<= x"20";
        when x"0BCC" => data_out<= x"29";
        when x"0BCD" => data_out<= x"AE";
        when x"0BCE" => data_out<= x"20";
        when x"0BCF" => data_out<= x"7B";
        when x"0BD0" => data_out<= x"B0";
        when x"0BD1" => data_out<= x"A0";
        when x"0BD2" => data_out<= x"05";
        when x"0BD3" => data_out<= x"20";
        when x"0BD4" => data_out<= x"4F";
        when x"0BD5" => data_out<= x"AF";
        when x"0BD6" => data_out<= x"85";
        when x"0BD7" => data_out<= x"14";
        when x"0BD8" => data_out<= x"86";
        when x"0BD9" => data_out<= x"15";
        when x"0BDA" => data_out<= x"A0";
        when x"0BDB" => data_out<= x"02";
        when x"0BDC" => data_out<= x"B1";
        when x"0BDD" => data_out<= x"0C";
        when x"0BDE" => data_out<= x"A8";
        when x"0BDF" => data_out<= x"B1";
        when x"0BE0" => data_out<= x"14";
        when x"0BE1" => data_out<= x"20";
        when x"0BE2" => data_out<= x"AF";
        when x"0BE3" => data_out<= x"8C";
        when x"0BE4" => data_out<= x"20";
        when x"0BE5" => data_out<= x"43";
        when x"0BE6" => data_out<= x"B0";
        when x"0BE7" => data_out<= x"A0";
        when x"0BE8" => data_out<= x"01";
        when x"0BE9" => data_out<= x"91";
        when x"0BEA" => data_out<= x"0C";
        when x"0BEB" => data_out<= x"88";
        when x"0BEC" => data_out<= x"B1";
        when x"0BED" => data_out<= x"0C";
        when x"0BEE" => data_out<= x"18";
        when x"0BEF" => data_out<= x"69";
        when x"0BF0" => data_out<= x"01";
        when x"0BF1" => data_out<= x"4C";
        when x"0BF2" => data_out<= x"97";
        when x"0BF3" => data_out<= x"8B";
        when x"0BF4" => data_out<= x"A0";
        when x"0BF5" => data_out<= x"01";
        when x"0BF6" => data_out<= x"A2";
        when x"0BF7" => data_out<= x"00";
        when x"0BF8" => data_out<= x"B1";
        when x"0BF9" => data_out<= x"0C";
        when x"0BFA" => data_out<= x"4C";
        when x"0BFB" => data_out<= x"27";
        when x"0BFC" => data_out<= x"AF";
        when x"0BFD" => data_out<= x"20";
        when x"0BFE" => data_out<= x"65";
        when x"0BFF" => data_out<= x"B0";
        when x"0C00" => data_out<= x"A0";
        when x"0C01" => data_out<= x"00";
        when x"0C02" => data_out<= x"B1";
        when x"0C03" => data_out<= x"0C";
        when x"0C04" => data_out<= x"4A";
        when x"0C05" => data_out<= x"4A";
        when x"0C06" => data_out<= x"4A";
        when x"0C07" => data_out<= x"4A";
        when x"0C08" => data_out<= x"29";
        when x"0C09" => data_out<= x"0F";
        when x"0C0A" => data_out<= x"85";
        when x"0C0B" => data_out<= x"14";
        when x"0C0C" => data_out<= x"98";
        when x"0C0D" => data_out<= x"18";
        when x"0C0E" => data_out<= x"69";
        when x"0C0F" => data_out<= x"B1";
        when x"0C10" => data_out<= x"85";
        when x"0C11" => data_out<= x"15";
        when x"0C12" => data_out<= x"A0";
        when x"0C13" => data_out<= x"D0";
        when x"0C14" => data_out<= x"B1";
        when x"0C15" => data_out<= x"14";
        when x"0C16" => data_out<= x"20";
        when x"0C17" => data_out<= x"F0";
        when x"0C18" => data_out<= x"80";
        when x"0C19" => data_out<= x"A0";
        when x"0C1A" => data_out<= x"00";
        when x"0C1B" => data_out<= x"B1";
        when x"0C1C" => data_out<= x"0C";
        when x"0C1D" => data_out<= x"29";
        when x"0C1E" => data_out<= x"0F";
        when x"0C1F" => data_out<= x"85";
        when x"0C20" => data_out<= x"14";
        when x"0C21" => data_out<= x"98";
        when x"0C22" => data_out<= x"18";
        when x"0C23" => data_out<= x"69";
        when x"0C24" => data_out<= x"B1";
        when x"0C25" => data_out<= x"85";
        when x"0C26" => data_out<= x"15";
        when x"0C27" => data_out<= x"A0";
        when x"0C28" => data_out<= x"D0";
        when x"0C29" => data_out<= x"B1";
        when x"0C2A" => data_out<= x"14";
        when x"0C2B" => data_out<= x"20";
        when x"0C2C" => data_out<= x"F0";
        when x"0C2D" => data_out<= x"80";
        when x"0C2E" => data_out<= x"4C";
        when x"0C2F" => data_out<= x"05";
        when x"0C30" => data_out<= x"AF";
        when x"0C31" => data_out<= x"20";
        when x"0C32" => data_out<= x"7B";
        when x"0C33" => data_out<= x"B0";
        when x"0C34" => data_out<= x"A0";
        when x"0C35" => data_out<= x"01";
        when x"0C36" => data_out<= x"B1";
        when x"0C37" => data_out<= x"0C";
        when x"0C38" => data_out<= x"20";
        when x"0C39" => data_out<= x"FD";
        when x"0C3A" => data_out<= x"8B";
        when x"0C3B" => data_out<= x"A0";
        when x"0C3C" => data_out<= x"00";
        when x"0C3D" => data_out<= x"B1";
        when x"0C3E" => data_out<= x"0C";
        when x"0C3F" => data_out<= x"20";
        when x"0C40" => data_out<= x"FD";
        when x"0C41" => data_out<= x"8B";
        when x"0C42" => data_out<= x"4C";
        when x"0C43" => data_out<= x"14";
        when x"0C44" => data_out<= x"AF";
        when x"0C45" => data_out<= x"A9";
        when x"0C46" => data_out<= x"0D";
        when x"0C47" => data_out<= x"20";
        when x"0C48" => data_out<= x"F0";
        when x"0C49" => data_out<= x"80";
        when x"0C4A" => data_out<= x"A9";
        when x"0C4B" => data_out<= x"0A";
        when x"0C4C" => data_out<= x"4C";
        when x"0C4D" => data_out<= x"F0";
        when x"0C4E" => data_out<= x"80";
        when x"0C4F" => data_out<= x"20";
        when x"0C50" => data_out<= x"7B";
        when x"0C51" => data_out<= x"B0";
        when x"0C52" => data_out<= x"20";
        when x"0C53" => data_out<= x"91";
        when x"0C54" => data_out<= x"B0";
        when x"0C55" => data_out<= x"A9";
        when x"0C56" => data_out<= x"D7";
        when x"0C57" => data_out<= x"A2";
        when x"0C58" => data_out<= x"BA";
        when x"0C59" => data_out<= x"20";
        when x"0C5A" => data_out<= x"22";
        when x"0C5B" => data_out<= x"81";
        when x"0C5C" => data_out<= x"A0";
        when x"0C5D" => data_out<= x"03";
        when x"0C5E" => data_out<= x"20";
        when x"0C5F" => data_out<= x"4F";
        when x"0C60" => data_out<= x"AF";
        when x"0C61" => data_out<= x"20";
        when x"0C62" => data_out<= x"31";
        when x"0C63" => data_out<= x"8C";
        when x"0C64" => data_out<= x"A9";
        when x"0C65" => data_out<= x"91";
        when x"0C66" => data_out<= x"A2";
        when x"0C67" => data_out<= x"B7";
        when x"0C68" => data_out<= x"20";
        when x"0C69" => data_out<= x"22";
        when x"0C6A" => data_out<= x"81";
        when x"0C6B" => data_out<= x"20";
        when x"0C6C" => data_out<= x"45";
        when x"0C6D" => data_out<= x"8C";
        when x"0C6E" => data_out<= x"20";
        when x"0C6F" => data_out<= x"4D";
        when x"0C70" => data_out<= x"AF";
        when x"0C71" => data_out<= x"20";
        when x"0C72" => data_out<= x"53";
        when x"0C73" => data_out<= x"AE";
        when x"0C74" => data_out<= x"20";
        when x"0C75" => data_out<= x"45";
        when x"0C76" => data_out<= x"8C";
        when x"0C77" => data_out<= x"A9";
        when x"0C78" => data_out<= x"97";
        when x"0C79" => data_out<= x"A2";
        when x"0C7A" => data_out<= x"BB";
        when x"0C7B" => data_out<= x"20";
        when x"0C7C" => data_out<= x"22";
        when x"0C7D" => data_out<= x"81";
        when x"0C7E" => data_out<= x"A0";
        when x"0C7F" => data_out<= x"03";
        when x"0C80" => data_out<= x"20";
        when x"0C81" => data_out<= x"4F";
        when x"0C82" => data_out<= x"AF";
        when x"0C83" => data_out<= x"20";
        when x"0C84" => data_out<= x"31";
        when x"0C85" => data_out<= x"8C";
        when x"0C86" => data_out<= x"20";
        when x"0C87" => data_out<= x"45";
        when x"0C88" => data_out<= x"8C";
        when x"0C89" => data_out<= x"4C";
        when x"0C8A" => data_out<= x"27";
        when x"0C8B" => data_out<= x"AF";
        when x"0C8C" => data_out<= x"A9";
        when x"0C8D" => data_out<= x"20";
        when x"0C8E" => data_out<= x"4C";
        when x"0C8F" => data_out<= x"F0";
        when x"0C90" => data_out<= x"80";
        when x"0C91" => data_out<= x"20";
        when x"0C92" => data_out<= x"45";
        when x"0C93" => data_out<= x"8C";
        when x"0C94" => data_out<= x"A9";
        when x"0C95" => data_out<= x"3E";
        when x"0C96" => data_out<= x"4C";
        when x"0C97" => data_out<= x"F0";
        when x"0C98" => data_out<= x"80";
        when x"0C99" => data_out<= x"20";
        when x"0C9A" => data_out<= x"7B";
        when x"0C9B" => data_out<= x"B0";
        when x"0C9C" => data_out<= x"A9";
        when x"0C9D" => data_out<= x"7F";
        when x"0C9E" => data_out<= x"A2";
        when x"0C9F" => data_out<= x"BC";
        when x"0CA0" => data_out<= x"20";
        when x"0CA1" => data_out<= x"22";
        when x"0CA2" => data_out<= x"81";
        when x"0CA3" => data_out<= x"20";
        when x"0CA4" => data_out<= x"4D";
        when x"0CA5" => data_out<= x"AF";
        when x"0CA6" => data_out<= x"20";
        when x"0CA7" => data_out<= x"22";
        when x"0CA8" => data_out<= x"81";
        when x"0CA9" => data_out<= x"20";
        when x"0CAA" => data_out<= x"45";
        when x"0CAB" => data_out<= x"8C";
        when x"0CAC" => data_out<= x"4C";
        when x"0CAD" => data_out<= x"14";
        when x"0CAE" => data_out<= x"AF";
        when x"0CAF" => data_out<= x"20";
        when x"0CB0" => data_out<= x"65";
        when x"0CB1" => data_out<= x"B0";
        when x"0CB2" => data_out<= x"A0";
        when x"0CB3" => data_out<= x"00";
        when x"0CB4" => data_out<= x"B1";
        when x"0CB5" => data_out<= x"0C";
        when x"0CB6" => data_out<= x"C9";
        when x"0CB7" => data_out<= x"30";
        when x"0CB8" => data_out<= x"90";
        when x"0CB9" => data_out<= x"12";
        when x"0CBA" => data_out<= x"C9";
        when x"0CBB" => data_out<= x"3A";
        when x"0CBC" => data_out<= x"B0";
        when x"0CBD" => data_out<= x"0E";
        when x"0CBE" => data_out<= x"A2";
        when x"0CBF" => data_out<= x"00";
        when x"0CC0" => data_out<= x"B1";
        when x"0CC1" => data_out<= x"0C";
        when x"0CC2" => data_out<= x"A0";
        when x"0CC3" => data_out<= x"30";
        when x"0CC4" => data_out<= x"20";
        when x"0CC5" => data_out<= x"61";
        when x"0CC6" => data_out<= x"AE";
        when x"0CC7" => data_out<= x"A2";
        when x"0CC8" => data_out<= x"00";
        when x"0CC9" => data_out<= x"4C";
        when x"0CCA" => data_out<= x"05";
        when x"0CCB" => data_out<= x"AF";
        when x"0CCC" => data_out<= x"B1";
        when x"0CCD" => data_out<= x"0C";
        when x"0CCE" => data_out<= x"C9";
        when x"0CCF" => data_out<= x"41";
        when x"0CD0" => data_out<= x"90";
        when x"0CD1" => data_out<= x"17";
        when x"0CD2" => data_out<= x"C9";
        when x"0CD3" => data_out<= x"47";
        when x"0CD4" => data_out<= x"B0";
        when x"0CD5" => data_out<= x"13";
        when x"0CD6" => data_out<= x"A2";
        when x"0CD7" => data_out<= x"00";
        when x"0CD8" => data_out<= x"B1";
        when x"0CD9" => data_out<= x"0C";
        when x"0CDA" => data_out<= x"A0";
        when x"0CDB" => data_out<= x"41";
        when x"0CDC" => data_out<= x"20";
        when x"0CDD" => data_out<= x"61";
        when x"0CDE" => data_out<= x"AE";
        when x"0CDF" => data_out<= x"A0";
        when x"0CE0" => data_out<= x"0A";
        when x"0CE1" => data_out<= x"20";
        when x"0CE2" => data_out<= x"FC";
        when x"0CE3" => data_out<= x"AE";
        when x"0CE4" => data_out<= x"A2";
        when x"0CE5" => data_out<= x"00";
        when x"0CE6" => data_out<= x"4C";
        when x"0CE7" => data_out<= x"05";
        when x"0CE8" => data_out<= x"AF";
        when x"0CE9" => data_out<= x"B1";
        when x"0CEA" => data_out<= x"0C";
        when x"0CEB" => data_out<= x"C9";
        when x"0CEC" => data_out<= x"61";
        when x"0CED" => data_out<= x"A2";
        when x"0CEE" => data_out<= x"00";
        when x"0CEF" => data_out<= x"90";
        when x"0CF0" => data_out<= x"15";
        when x"0CF1" => data_out<= x"B1";
        when x"0CF2" => data_out<= x"0C";
        when x"0CF3" => data_out<= x"C9";
        when x"0CF4" => data_out<= x"67";
        when x"0CF5" => data_out<= x"B0";
        when x"0CF6" => data_out<= x"0F";
        when x"0CF7" => data_out<= x"A0";
        when x"0CF8" => data_out<= x"61";
        when x"0CF9" => data_out<= x"20";
        when x"0CFA" => data_out<= x"61";
        when x"0CFB" => data_out<= x"AE";
        when x"0CFC" => data_out<= x"A0";
        when x"0CFD" => data_out<= x"0A";
        when x"0CFE" => data_out<= x"20";
        when x"0CFF" => data_out<= x"FC";
        when x"0D00" => data_out<= x"AE";
        when x"0D01" => data_out<= x"A2";
        when x"0D02" => data_out<= x"00";
        when x"0D03" => data_out<= x"4C";
        when x"0D04" => data_out<= x"05";
        when x"0D05" => data_out<= x"AF";
        when x"0D06" => data_out<= x"A9";
        when x"0D07" => data_out<= x"FF";
        when x"0D08" => data_out<= x"4C";
        when x"0D09" => data_out<= x"05";
        when x"0D0A" => data_out<= x"AF";
        when x"0D0B" => data_out<= x"20";
        when x"0D0C" => data_out<= x"65";
        when x"0D0D" => data_out<= x"B0";
        when x"0D0E" => data_out<= x"A0";
        when x"0D0F" => data_out<= x"00";
        when x"0D10" => data_out<= x"B1";
        when x"0D11" => data_out<= x"0C";
        when x"0D12" => data_out<= x"C9";
        when x"0D13" => data_out<= x"30";
        when x"0D14" => data_out<= x"90";
        when x"0D15" => data_out<= x"0D";
        when x"0D16" => data_out<= x"A2";
        when x"0D17" => data_out<= x"00";
        when x"0D18" => data_out<= x"B1";
        when x"0D19" => data_out<= x"0C";
        when x"0D1A" => data_out<= x"C9";
        when x"0D1B" => data_out<= x"3A";
        when x"0D1C" => data_out<= x"B0";
        when x"0D1D" => data_out<= x"05";
        when x"0D1E" => data_out<= x"A9";
        when x"0D1F" => data_out<= x"01";
        when x"0D20" => data_out<= x"4C";
        when x"0D21" => data_out<= x"05";
        when x"0D22" => data_out<= x"AF";
        when x"0D23" => data_out<= x"B1";
        when x"0D24" => data_out<= x"0C";
        when x"0D25" => data_out<= x"C9";
        when x"0D26" => data_out<= x"41";
        when x"0D27" => data_out<= x"90";
        when x"0D28" => data_out<= x"0D";
        when x"0D29" => data_out<= x"A2";
        when x"0D2A" => data_out<= x"00";
        when x"0D2B" => data_out<= x"B1";
        when x"0D2C" => data_out<= x"0C";
        when x"0D2D" => data_out<= x"C9";
        when x"0D2E" => data_out<= x"47";
        when x"0D2F" => data_out<= x"B0";
        when x"0D30" => data_out<= x"05";
        when x"0D31" => data_out<= x"A9";
        when x"0D32" => data_out<= x"01";
        when x"0D33" => data_out<= x"4C";
        when x"0D34" => data_out<= x"05";
        when x"0D35" => data_out<= x"AF";
        when x"0D36" => data_out<= x"B1";
        when x"0D37" => data_out<= x"0C";
        when x"0D38" => data_out<= x"C9";
        when x"0D39" => data_out<= x"61";
        when x"0D3A" => data_out<= x"98";
        when x"0D3B" => data_out<= x"AA";
        when x"0D3C" => data_out<= x"90";
        when x"0D3D" => data_out<= x"0F";
        when x"0D3E" => data_out<= x"B1";
        when x"0D3F" => data_out<= x"0C";
        when x"0D40" => data_out<= x"C9";
        when x"0D41" => data_out<= x"67";
        when x"0D42" => data_out<= x"90";
        when x"0D43" => data_out<= x"04";
        when x"0D44" => data_out<= x"8A";
        when x"0D45" => data_out<= x"4C";
        when x"0D46" => data_out<= x"05";
        when x"0D47" => data_out<= x"AF";
        when x"0D48" => data_out<= x"A9";
        when x"0D49" => data_out<= x"01";
        when x"0D4A" => data_out<= x"4C";
        when x"0D4B" => data_out<= x"05";
        when x"0D4C" => data_out<= x"AF";
        when x"0D4D" => data_out<= x"4C";
        when x"0D4E" => data_out<= x"05";
        when x"0D4F" => data_out<= x"AF";
        when x"0D50" => data_out<= x"20";
        when x"0D51" => data_out<= x"7B";
        when x"0D52" => data_out<= x"B0";
        when x"0D53" => data_out<= x"20";
        when x"0D54" => data_out<= x"4D";
        when x"0D55" => data_out<= x"AF";
        when x"0D56" => data_out<= x"85";
        when x"0D57" => data_out<= x"14";
        when x"0D58" => data_out<= x"86";
        when x"0D59" => data_out<= x"15";
        when x"0D5A" => data_out<= x"A9";
        when x"0D5B" => data_out<= x"00";
        when x"0D5C" => data_out<= x"A8";
        when x"0D5D" => data_out<= x"91";
        when x"0D5E" => data_out<= x"14";
        when x"0D5F" => data_out<= x"C8";
        when x"0D60" => data_out<= x"91";
        when x"0D61" => data_out<= x"14";
        when x"0D62" => data_out<= x"4C";
        when x"0D63" => data_out<= x"72";
        when x"0D64" => data_out<= x"8D";
        when x"0D65" => data_out<= x"A0";
        when x"0D66" => data_out<= x"03";
        when x"0D67" => data_out<= x"20";
        when x"0D68" => data_out<= x"4F";
        when x"0D69" => data_out<= x"AF";
        when x"0D6A" => data_out<= x"20";
        when x"0D6B" => data_out<= x"E2";
        when x"0D6C" => data_out<= x"AE";
        when x"0D6D" => data_out<= x"A0";
        when x"0D6E" => data_out<= x"02";
        when x"0D6F" => data_out<= x"20";
        when x"0D70" => data_out<= x"C5";
        when x"0D71" => data_out<= x"B0";
        when x"0D72" => data_out<= x"A0";
        when x"0D73" => data_out<= x"03";
        when x"0D74" => data_out<= x"20";
        when x"0D75" => data_out<= x"4F";
        when x"0D76" => data_out<= x"AF";
        when x"0D77" => data_out<= x"85";
        when x"0D78" => data_out<= x"14";
        when x"0D79" => data_out<= x"86";
        when x"0D7A" => data_out<= x"15";
        when x"0D7B" => data_out<= x"A0";
        when x"0D7C" => data_out<= x"00";
        when x"0D7D" => data_out<= x"B1";
        when x"0D7E" => data_out<= x"14";
        when x"0D7F" => data_out<= x"C9";
        when x"0D80" => data_out<= x"20";
        when x"0D81" => data_out<= x"F0";
        when x"0D82" => data_out<= x"E2";
        when x"0D83" => data_out<= x"4C";
        when x"0D84" => data_out<= x"BC";
        when x"0D85" => data_out<= x"8D";
        when x"0D86" => data_out<= x"20";
        when x"0D87" => data_out<= x"91";
        when x"0D88" => data_out<= x"B0";
        when x"0D89" => data_out<= x"A0";
        when x"0D8A" => data_out<= x"03";
        when x"0D8B" => data_out<= x"20";
        when x"0D8C" => data_out<= x"4F";
        when x"0D8D" => data_out<= x"AF";
        when x"0D8E" => data_out<= x"20";
        when x"0D8F" => data_out<= x"40";
        when x"0D90" => data_out<= x"AF";
        when x"0D91" => data_out<= x"20";
        when x"0D92" => data_out<= x"29";
        when x"0D93" => data_out<= x"AE";
        when x"0D94" => data_out<= x"20";
        when x"0D95" => data_out<= x"7B";
        when x"0D96" => data_out<= x"B0";
        when x"0D97" => data_out<= x"A0";
        when x"0D98" => data_out<= x"07";
        when x"0D99" => data_out<= x"20";
        when x"0D9A" => data_out<= x"4F";
        when x"0D9B" => data_out<= x"AF";
        when x"0D9C" => data_out<= x"85";
        when x"0D9D" => data_out<= x"14";
        when x"0D9E" => data_out<= x"86";
        when x"0D9F" => data_out<= x"15";
        when x"0DA0" => data_out<= x"A0";
        when x"0DA1" => data_out<= x"00";
        when x"0DA2" => data_out<= x"B1";
        when x"0DA3" => data_out<= x"14";
        when x"0DA4" => data_out<= x"20";
        when x"0DA5" => data_out<= x"AF";
        when x"0DA6" => data_out<= x"8C";
        when x"0DA7" => data_out<= x"20";
        when x"0DA8" => data_out<= x"43";
        when x"0DA9" => data_out<= x"B0";
        when x"0DAA" => data_out<= x"A0";
        when x"0DAB" => data_out<= x"00";
        when x"0DAC" => data_out<= x"20";
        when x"0DAD" => data_out<= x"CE";
        when x"0DAE" => data_out<= x"B0";
        when x"0DAF" => data_out<= x"A0";
        when x"0DB0" => data_out<= x"03";
        when x"0DB1" => data_out<= x"20";
        when x"0DB2" => data_out<= x"4F";
        when x"0DB3" => data_out<= x"AF";
        when x"0DB4" => data_out<= x"20";
        when x"0DB5" => data_out<= x"E2";
        when x"0DB6" => data_out<= x"AE";
        when x"0DB7" => data_out<= x"A0";
        when x"0DB8" => data_out<= x"02";
        when x"0DB9" => data_out<= x"20";
        when x"0DBA" => data_out<= x"C5";
        when x"0DBB" => data_out<= x"B0";
        when x"0DBC" => data_out<= x"A0";
        when x"0DBD" => data_out<= x"03";
        when x"0DBE" => data_out<= x"20";
        when x"0DBF" => data_out<= x"4F";
        when x"0DC0" => data_out<= x"AF";
        when x"0DC1" => data_out<= x"85";
        when x"0DC2" => data_out<= x"14";
        when x"0DC3" => data_out<= x"86";
        when x"0DC4" => data_out<= x"15";
        when x"0DC5" => data_out<= x"A0";
        when x"0DC6" => data_out<= x"00";
        when x"0DC7" => data_out<= x"B1";
        when x"0DC8" => data_out<= x"14";
        when x"0DC9" => data_out<= x"20";
        when x"0DCA" => data_out<= x"0B";
        when x"0DCB" => data_out<= x"8D";
        when x"0DCC" => data_out<= x"AA";
        when x"0DCD" => data_out<= x"D0";
        when x"0DCE" => data_out<= x"B7";
        when x"0DCF" => data_out<= x"A0";
        when x"0DD0" => data_out<= x"03";
        when x"0DD1" => data_out<= x"20";
        when x"0DD2" => data_out<= x"4F";
        when x"0DD3" => data_out<= x"AF";
        when x"0DD4" => data_out<= x"4C";
        when x"0DD5" => data_out<= x"27";
        when x"0DD6" => data_out<= x"AF";
        when x"0DD7" => data_out<= x"20";
        when x"0DD8" => data_out<= x"7B";
        when x"0DD9" => data_out<= x"B0";
        when x"0DDA" => data_out<= x"20";
        when x"0DDB" => data_out<= x"73";
        when x"0DDC" => data_out<= x"AE";
        when x"0DDD" => data_out<= x"A9";
        when x"0DDE" => data_out<= x"00";
        when x"0DDF" => data_out<= x"20";
        when x"0DE0" => data_out<= x"65";
        when x"0DE1" => data_out<= x"B0";
        when x"0DE2" => data_out<= x"20";
        when x"0DE3" => data_out<= x"77";
        when x"0DE4" => data_out<= x"B0";
        when x"0DE5" => data_out<= x"A9";
        when x"0DE6" => data_out<= x"17";
        when x"0DE7" => data_out<= x"A2";
        when x"0DE8" => data_out<= x"BB";
        when x"0DE9" => data_out<= x"20";
        when x"0DEA" => data_out<= x"22";
        when x"0DEB" => data_out<= x"81";
        when x"0DEC" => data_out<= x"A0";
        when x"0DED" => data_out<= x"06";
        when x"0DEE" => data_out<= x"20";
        when x"0DEF" => data_out<= x"4F";
        when x"0DF0" => data_out<= x"AF";
        when x"0DF1" => data_out<= x"20";
        when x"0DF2" => data_out<= x"31";
        when x"0DF3" => data_out<= x"8C";
        when x"0DF4" => data_out<= x"A9";
        when x"0DF5" => data_out<= x"D4";
        when x"0DF6" => data_out<= x"A2";
        when x"0DF7" => data_out<= x"B9";
        when x"0DF8" => data_out<= x"20";
        when x"0DF9" => data_out<= x"22";
        when x"0DFA" => data_out<= x"81";
        when x"0DFB" => data_out<= x"20";
        when x"0DFC" => data_out<= x"45";
        when x"0DFD" => data_out<= x"8C";
        when x"0DFE" => data_out<= x"A9";
        when x"0DFF" => data_out<= x"3A";
        when x"0E00" => data_out<= x"20";
        when x"0E01" => data_out<= x"F0";
        when x"0E02" => data_out<= x"80";
        when x"0E03" => data_out<= x"A9";
        when x"0E04" => data_out<= x"00";
        when x"0E05" => data_out<= x"A0";
        when x"0E06" => data_out<= x"03";
        when x"0E07" => data_out<= x"91";
        when x"0E08" => data_out<= x"0C";
        when x"0E09" => data_out<= x"20";
        when x"0E0A" => data_out<= x"FD";
        when x"0E0B" => data_out<= x"80";
        when x"0E0C" => data_out<= x"A0";
        when x"0E0D" => data_out<= x"04";
        when x"0E0E" => data_out<= x"91";
        when x"0E0F" => data_out<= x"0C";
        when x"0E10" => data_out<= x"C9";
        when x"0E11" => data_out<= x"2E";
        when x"0E12" => data_out<= x"D0";
        when x"0E13" => data_out<= x"03";
        when x"0E14" => data_out<= x"4C";
        when x"0E15" => data_out<= x"99";
        when x"0E16" => data_out<= x"8E";
        when x"0E17" => data_out<= x"B1";
        when x"0E18" => data_out<= x"0C";
        when x"0E19" => data_out<= x"C9";
        when x"0E1A" => data_out<= x"0D";
        when x"0E1B" => data_out<= x"F0";
        when x"0E1C" => data_out<= x"04";
        when x"0E1D" => data_out<= x"C9";
        when x"0E1E" => data_out<= x"0A";
        when x"0E1F" => data_out<= x"D0";
        when x"0E20" => data_out<= x"0B";
        when x"0E21" => data_out<= x"20";
        when x"0E22" => data_out<= x"45";
        when x"0E23" => data_out<= x"8C";
        when x"0E24" => data_out<= x"A9";
        when x"0E25" => data_out<= x"3A";
        when x"0E26" => data_out<= x"20";
        when x"0E27" => data_out<= x"F0";
        when x"0E28" => data_out<= x"80";
        when x"0E29" => data_out<= x"4C";
        when x"0E2A" => data_out<= x"09";
        when x"0E2B" => data_out<= x"8E";
        when x"0E2C" => data_out<= x"B1";
        when x"0E2D" => data_out<= x"0C";
        when x"0E2E" => data_out<= x"C9";
        when x"0E2F" => data_out<= x"20";
        when x"0E30" => data_out<= x"D0";
        when x"0E31" => data_out<= x"06";
        when x"0E32" => data_out<= x"20";
        when x"0E33" => data_out<= x"F0";
        when x"0E34" => data_out<= x"80";
        when x"0E35" => data_out<= x"4C";
        when x"0E36" => data_out<= x"09";
        when x"0E37" => data_out<= x"8E";
        when x"0E38" => data_out<= x"B1";
        when x"0E39" => data_out<= x"0C";
        when x"0E3A" => data_out<= x"20";
        when x"0E3B" => data_out<= x"0B";
        when x"0E3C" => data_out<= x"8D";
        when x"0E3D" => data_out<= x"AA";
        when x"0E3E" => data_out<= x"F0";
        when x"0E3F" => data_out<= x"C9";
        when x"0E40" => data_out<= x"A0";
        when x"0E41" => data_out<= x"04";
        when x"0E42" => data_out<= x"B1";
        when x"0E43" => data_out<= x"0C";
        when x"0E44" => data_out<= x"20";
        when x"0E45" => data_out<= x"F0";
        when x"0E46" => data_out<= x"80";
        when x"0E47" => data_out<= x"A0";
        when x"0E48" => data_out<= x"03";
        when x"0E49" => data_out<= x"A2";
        when x"0E4A" => data_out<= x"00";
        when x"0E4B" => data_out<= x"B1";
        when x"0E4C" => data_out<= x"0C";
        when x"0E4D" => data_out<= x"20";
        when x"0E4E" => data_out<= x"29";
        when x"0E4F" => data_out<= x"AE";
        when x"0E50" => data_out<= x"20";
        when x"0E51" => data_out<= x"7B";
        when x"0E52" => data_out<= x"B0";
        when x"0E53" => data_out<= x"A0";
        when x"0E54" => data_out<= x"06";
        when x"0E55" => data_out<= x"B1";
        when x"0E56" => data_out<= x"0C";
        when x"0E57" => data_out<= x"20";
        when x"0E58" => data_out<= x"AF";
        when x"0E59" => data_out<= x"8C";
        when x"0E5A" => data_out<= x"20";
        when x"0E5B" => data_out<= x"43";
        when x"0E5C" => data_out<= x"B0";
        when x"0E5D" => data_out<= x"A0";
        when x"0E5E" => data_out<= x"03";
        when x"0E5F" => data_out<= x"91";
        when x"0E60" => data_out<= x"0C";
        when x"0E61" => data_out<= x"88";
        when x"0E62" => data_out<= x"B1";
        when x"0E63" => data_out<= x"0C";
        when x"0E64" => data_out<= x"18";
        when x"0E65" => data_out<= x"69";
        when x"0E66" => data_out<= x"01";
        when x"0E67" => data_out<= x"91";
        when x"0E68" => data_out<= x"0C";
        when x"0E69" => data_out<= x"C9";
        when x"0E6A" => data_out<= x"02";
        when x"0E6B" => data_out<= x"D0";
        when x"0E6C" => data_out<= x"9C";
        when x"0E6D" => data_out<= x"A0";
        when x"0E6E" => data_out<= x"08";
        when x"0E6F" => data_out<= x"20";
        when x"0E70" => data_out<= x"93";
        when x"0E71" => data_out<= x"B0";
        when x"0E72" => data_out<= x"A0";
        when x"0E73" => data_out<= x"05";
        when x"0E74" => data_out<= x"B1";
        when x"0E75" => data_out<= x"0C";
        when x"0E76" => data_out<= x"20";
        when x"0E77" => data_out<= x"5A";
        when x"0E78" => data_out<= x"89";
        when x"0E79" => data_out<= x"A0";
        when x"0E7A" => data_out<= x"06";
        when x"0E7B" => data_out<= x"20";
        when x"0E7C" => data_out<= x"4F";
        when x"0E7D" => data_out<= x"AF";
        when x"0E7E" => data_out<= x"20";
        when x"0E7F" => data_out<= x"E2";
        when x"0E80" => data_out<= x"AE";
        when x"0E81" => data_out<= x"A0";
        when x"0E82" => data_out<= x"05";
        when x"0E83" => data_out<= x"20";
        when x"0E84" => data_out<= x"C5";
        when x"0E85" => data_out<= x"B0";
        when x"0E86" => data_out<= x"20";
        when x"0E87" => data_out<= x"4D";
        when x"0E88" => data_out<= x"AF";
        when x"0E89" => data_out<= x"20";
        when x"0E8A" => data_out<= x"E2";
        when x"0E8B" => data_out<= x"AE";
        when x"0E8C" => data_out<= x"20";
        when x"0E8D" => data_out<= x"C3";
        when x"0E8E" => data_out<= x"B0";
        when x"0E8F" => data_out<= x"A9";
        when x"0E90" => data_out<= x"00";
        when x"0E91" => data_out<= x"A0";
        when x"0E92" => data_out<= x"03";
        when x"0E93" => data_out<= x"91";
        when x"0E94" => data_out<= x"0C";
        when x"0E95" => data_out<= x"88";
        when x"0E96" => data_out<= x"4C";
        when x"0E97" => data_out<= x"07";
        when x"0E98" => data_out<= x"8E";
        when x"0E99" => data_out<= x"20";
        when x"0E9A" => data_out<= x"45";
        when x"0E9B" => data_out<= x"8C";
        when x"0E9C" => data_out<= x"A9";
        when x"0E9D" => data_out<= x"E2";
        when x"0E9E" => data_out<= x"A2";
        when x"0E9F" => data_out<= x"BB";
        when x"0EA0" => data_out<= x"20";
        when x"0EA1" => data_out<= x"22";
        when x"0EA2" => data_out<= x"81";
        when x"0EA3" => data_out<= x"20";
        when x"0EA4" => data_out<= x"4D";
        when x"0EA5" => data_out<= x"AF";
        when x"0EA6" => data_out<= x"20";
        when x"0EA7" => data_out<= x"31";
        when x"0EA8" => data_out<= x"8C";
        when x"0EA9" => data_out<= x"A9";
        when x"0EAA" => data_out<= x"34";
        when x"0EAB" => data_out<= x"A2";
        when x"0EAC" => data_out<= x"BC";
        when x"0EAD" => data_out<= x"20";
        when x"0EAE" => data_out<= x"22";
        when x"0EAF" => data_out<= x"81";
        when x"0EB0" => data_out<= x"20";
        when x"0EB1" => data_out<= x"45";
        when x"0EB2" => data_out<= x"8C";
        when x"0EB3" => data_out<= x"A0";
        when x"0EB4" => data_out<= x"06";
        when x"0EB5" => data_out<= x"20";
        when x"0EB6" => data_out<= x"4F";
        when x"0EB7" => data_out<= x"AF";
        when x"0EB8" => data_out<= x"8D";
        when x"0EB9" => data_out<= x"00";
        when x"0EBA" => data_out<= x"02";
        when x"0EBB" => data_out<= x"8E";
        when x"0EBC" => data_out<= x"01";
        when x"0EBD" => data_out<= x"02";
        when x"0EBE" => data_out<= x"4C";
        when x"0EBF" => data_out<= x"36";
        when x"0EC0" => data_out<= x"AF";
        when x"0EC1" => data_out<= x"20";
        when x"0EC2" => data_out<= x"65";
        when x"0EC3" => data_out<= x"B0";
        when x"0EC4" => data_out<= x"A0";
        when x"0EC5" => data_out<= x"00";
        when x"0EC6" => data_out<= x"B1";
        when x"0EC7" => data_out<= x"0C";
        when x"0EC8" => data_out<= x"D0";
        when x"0EC9" => data_out<= x"03";
        when x"0ECA" => data_out<= x"4C";
        when x"0ECB" => data_out<= x"35";
        when x"0ECC" => data_out<= x"90";
        when x"0ECD" => data_out<= x"C9";
        when x"0ECE" => data_out<= x"08";
        when x"0ECF" => data_out<= x"D0";
        when x"0ED0" => data_out<= x"03";
        when x"0ED1" => data_out<= x"4C";
        when x"0ED2" => data_out<= x"23";
        when x"0ED3" => data_out<= x"91";
        when x"0ED4" => data_out<= x"C9";
        when x"0ED5" => data_out<= x"09";
        when x"0ED6" => data_out<= x"D0";
        when x"0ED7" => data_out<= x"03";
        when x"0ED8" => data_out<= x"4C";
        when x"0ED9" => data_out<= x"5B";
        when x"0EDA" => data_out<= x"91";
        when x"0EDB" => data_out<= x"C9";
        when x"0EDC" => data_out<= x"10";
        when x"0EDD" => data_out<= x"D0";
        when x"0EDE" => data_out<= x"03";
        when x"0EDF" => data_out<= x"4C";
        when x"0EE0" => data_out<= x"77";
        when x"0EE1" => data_out<= x"91";
        when x"0EE2" => data_out<= x"C9";
        when x"0EE3" => data_out<= x"18";
        when x"0EE4" => data_out<= x"D0";
        when x"0EE5" => data_out<= x"03";
        when x"0EE6" => data_out<= x"4C";
        when x"0EE7" => data_out<= x"BA";
        when x"0EE8" => data_out<= x"90";
        when x"0EE9" => data_out<= x"C9";
        when x"0EEA" => data_out<= x"20";
        when x"0EEB" => data_out<= x"D0";
        when x"0EEC" => data_out<= x"03";
        when x"0EED" => data_out<= x"4C";
        when x"0EEE" => data_out<= x"3C";
        when x"0EEF" => data_out<= x"90";
        when x"0EF0" => data_out<= x"C9";
        when x"0EF1" => data_out<= x"28";
        when x"0EF2" => data_out<= x"D0";
        when x"0EF3" => data_out<= x"03";
        when x"0EF4" => data_out<= x"4C";
        when x"0EF5" => data_out<= x"2A";
        when x"0EF6" => data_out<= x"91";
        when x"0EF7" => data_out<= x"C9";
        when x"0EF8" => data_out<= x"29";
        when x"0EF9" => data_out<= x"D0";
        when x"0EFA" => data_out<= x"03";
        when x"0EFB" => data_out<= x"4C";
        when x"0EFC" => data_out<= x"54";
        when x"0EFD" => data_out<= x"91";
        when x"0EFE" => data_out<= x"C9";
        when x"0EFF" => data_out<= x"30";
        when x"0F00" => data_out<= x"D0";
        when x"0F01" => data_out<= x"03";
        when x"0F02" => data_out<= x"4C";
        when x"0F03" => data_out<= x"7E";
        when x"0F04" => data_out<= x"91";
        when x"0F05" => data_out<= x"C9";
        when x"0F06" => data_out<= x"38";
        when x"0F07" => data_out<= x"D0";
        when x"0F08" => data_out<= x"03";
        when x"0F09" => data_out<= x"4C";
        when x"0F0A" => data_out<= x"C1";
        when x"0F0B" => data_out<= x"90";
        when x"0F0C" => data_out<= x"C9";
        when x"0F0D" => data_out<= x"40";
        when x"0F0E" => data_out<= x"D0";
        when x"0F0F" => data_out<= x"03";
        when x"0F10" => data_out<= x"4C";
        when x"0F11" => data_out<= x"43";
        when x"0F12" => data_out<= x"90";
        when x"0F13" => data_out<= x"C9";
        when x"0F14" => data_out<= x"48";
        when x"0F15" => data_out<= x"D0";
        when x"0F16" => data_out<= x"03";
        when x"0F17" => data_out<= x"4C";
        when x"0F18" => data_out<= x"15";
        when x"0F19" => data_out<= x"91";
        when x"0F1A" => data_out<= x"C9";
        when x"0F1B" => data_out<= x"49";
        when x"0F1C" => data_out<= x"D0";
        when x"0F1D" => data_out<= x"03";
        when x"0F1E" => data_out<= x"4C";
        when x"0F1F" => data_out<= x"62";
        when x"0F20" => data_out<= x"91";
        when x"0F21" => data_out<= x"C9";
        when x"0F22" => data_out<= x"4C";
        when x"0F23" => data_out<= x"D0";
        when x"0F24" => data_out<= x"03";
        when x"0F25" => data_out<= x"4C";
        when x"0F26" => data_out<= x"51";
        when x"0F27" => data_out<= x"90";
        when x"0F28" => data_out<= x"C9";
        when x"0F29" => data_out<= x"50";
        when x"0F2A" => data_out<= x"D0";
        when x"0F2B" => data_out<= x"03";
        when x"0F2C" => data_out<= x"4C";
        when x"0F2D" => data_out<= x"93";
        when x"0F2E" => data_out<= x"91";
        when x"0F2F" => data_out<= x"C9";
        when x"0F30" => data_out<= x"58";
        when x"0F31" => data_out<= x"D0";
        when x"0F32" => data_out<= x"03";
        when x"0F33" => data_out<= x"4C";
        when x"0F34" => data_out<= x"D6";
        when x"0F35" => data_out<= x"90";
        when x"0F36" => data_out<= x"C9";
        when x"0F37" => data_out<= x"60";
        when x"0F38" => data_out<= x"D0";
        when x"0F39" => data_out<= x"03";
        when x"0F3A" => data_out<= x"4C";
        when x"0F3B" => data_out<= x"4A";
        when x"0F3C" => data_out<= x"90";
        when x"0F3D" => data_out<= x"C9";
        when x"0F3E" => data_out<= x"68";
        when x"0F3F" => data_out<= x"D0";
        when x"0F40" => data_out<= x"03";
        when x"0F41" => data_out<= x"4C";
        when x"0F42" => data_out<= x"1C";
        when x"0F43" => data_out<= x"91";
        when x"0F44" => data_out<= x"C9";
        when x"0F45" => data_out<= x"69";
        when x"0F46" => data_out<= x"D0";
        when x"0F47" => data_out<= x"03";
        when x"0F48" => data_out<= x"4C";
        when x"0F49" => data_out<= x"31";
        when x"0F4A" => data_out<= x"91";
        when x"0F4B" => data_out<= x"C9";
        when x"0F4C" => data_out<= x"6C";
        when x"0F4D" => data_out<= x"D0";
        when x"0F4E" => data_out<= x"03";
        when x"0F4F" => data_out<= x"4C";
        when x"0F50" => data_out<= x"58";
        when x"0F51" => data_out<= x"90";
        when x"0F52" => data_out<= x"C9";
        when x"0F53" => data_out<= x"70";
        when x"0F54" => data_out<= x"D0";
        when x"0F55" => data_out<= x"03";
        when x"0F56" => data_out<= x"4C";
        when x"0F57" => data_out<= x"9A";
        when x"0F58" => data_out<= x"91";
        when x"0F59" => data_out<= x"C9";
        when x"0F5A" => data_out<= x"78";
        when x"0F5B" => data_out<= x"D0";
        when x"0F5C" => data_out<= x"03";
        when x"0F5D" => data_out<= x"4C";
        when x"0F5E" => data_out<= x"DD";
        when x"0F5F" => data_out<= x"90";
        when x"0F60" => data_out<= x"C9";
        when x"0F61" => data_out<= x"84";
        when x"0F62" => data_out<= x"D0";
        when x"0F63" => data_out<= x"03";
        when x"0F64" => data_out<= x"4C";
        when x"0F65" => data_out<= x"97";
        when x"0F66" => data_out<= x"90";
        when x"0F67" => data_out<= x"C9";
        when x"0F68" => data_out<= x"85";
        when x"0F69" => data_out<= x"D0";
        when x"0F6A" => data_out<= x"03";
        when x"0F6B" => data_out<= x"4C";
        when x"0F6C" => data_out<= x"82";
        when x"0F6D" => data_out<= x"90";
        when x"0F6E" => data_out<= x"C9";
        when x"0F6F" => data_out<= x"86";
        when x"0F70" => data_out<= x"D0";
        when x"0F71" => data_out<= x"03";
        when x"0F72" => data_out<= x"4C";
        when x"0F73" => data_out<= x"90";
        when x"0F74" => data_out<= x"90";
        when x"0F75" => data_out<= x"C9";
        when x"0F76" => data_out<= x"88";
        when x"0F77" => data_out<= x"D0";
        when x"0F78" => data_out<= x"03";
        when x"0F79" => data_out<= x"4C";
        when x"0F7A" => data_out<= x"B3";
        when x"0F7B" => data_out<= x"90";
        when x"0F7C" => data_out<= x"C9";
        when x"0F7D" => data_out<= x"8A";
        when x"0F7E" => data_out<= x"D0";
        when x"0F7F" => data_out<= x"03";
        when x"0F80" => data_out<= x"4C";
        when x"0F81" => data_out<= x"F9";
        when x"0F82" => data_out<= x"90";
        when x"0F83" => data_out<= x"C9";
        when x"0F84" => data_out<= x"8D";
        when x"0F85" => data_out<= x"D0";
        when x"0F86" => data_out<= x"03";
        when x"0F87" => data_out<= x"4C";
        when x"0F88" => data_out<= x"89";
        when x"0F89" => data_out<= x"90";
        when x"0F8A" => data_out<= x"C9";
        when x"0F8B" => data_out<= x"90";
        when x"0F8C" => data_out<= x"D0";
        when x"0F8D" => data_out<= x"03";
        when x"0F8E" => data_out<= x"4C";
        when x"0F8F" => data_out<= x"85";
        when x"0F90" => data_out<= x"91";
        when x"0F91" => data_out<= x"C9";
        when x"0F92" => data_out<= x"98";
        when x"0F93" => data_out<= x"D0";
        when x"0F94" => data_out<= x"03";
        when x"0F95" => data_out<= x"4C";
        when x"0F96" => data_out<= x"00";
        when x"0F97" => data_out<= x"91";
        when x"0F98" => data_out<= x"C9";
        when x"0F99" => data_out<= x"9A";
        when x"0F9A" => data_out<= x"D0";
        when x"0F9B" => data_out<= x"03";
        when x"0F9C" => data_out<= x"4C";
        when x"0F9D" => data_out<= x"07";
        when x"0F9E" => data_out<= x"91";
        when x"0F9F" => data_out<= x"C9";
        when x"0FA0" => data_out<= x"A0";
        when x"0FA1" => data_out<= x"D0";
        when x"0FA2" => data_out<= x"03";
        when x"0FA3" => data_out<= x"4C";
        when x"0FA4" => data_out<= x"7B";
        when x"0FA5" => data_out<= x"90";
        when x"0FA6" => data_out<= x"C9";
        when x"0FA7" => data_out<= x"A2";
        when x"0FA8" => data_out<= x"D0";
        when x"0FA9" => data_out<= x"03";
        when x"0FAA" => data_out<= x"4C";
        when x"0FAB" => data_out<= x"74";
        when x"0FAC" => data_out<= x"90";
        when x"0FAD" => data_out<= x"C9";
        when x"0FAE" => data_out<= x"A5";
        when x"0FAF" => data_out<= x"D0";
        when x"0FB0" => data_out<= x"03";
        when x"0FB1" => data_out<= x"4C";
        when x"0FB2" => data_out<= x"66";
        when x"0FB3" => data_out<= x"90";
        when x"0FB4" => data_out<= x"C9";
        when x"0FB5" => data_out<= x"A8";
        when x"0FB6" => data_out<= x"D0";
        when x"0FB7" => data_out<= x"03";
        when x"0FB8" => data_out<= x"4C";
        when x"0FB9" => data_out<= x"F2";
        when x"0FBA" => data_out<= x"90";
        when x"0FBB" => data_out<= x"C9";
        when x"0FBC" => data_out<= x"A9";
        when x"0FBD" => data_out<= x"D0";
        when x"0FBE" => data_out<= x"03";
        when x"0FBF" => data_out<= x"4C";
        when x"0FC0" => data_out<= x"5F";
        when x"0FC1" => data_out<= x"90";
        when x"0FC2" => data_out<= x"C9";
        when x"0FC3" => data_out<= x"AA";
        when x"0FC4" => data_out<= x"D0";
        when x"0FC5" => data_out<= x"03";
        when x"0FC6" => data_out<= x"4C";
        when x"0FC7" => data_out<= x"EB";
        when x"0FC8" => data_out<= x"90";
        when x"0FC9" => data_out<= x"C9";
        when x"0FCA" => data_out<= x"AD";
        when x"0FCB" => data_out<= x"D0";
        when x"0FCC" => data_out<= x"03";
        when x"0FCD" => data_out<= x"4C";
        when x"0FCE" => data_out<= x"6D";
        when x"0FCF" => data_out<= x"90";
        when x"0FD0" => data_out<= x"C9";
        when x"0FD1" => data_out<= x"B0";
        when x"0FD2" => data_out<= x"D0";
        when x"0FD3" => data_out<= x"03";
        when x"0FD4" => data_out<= x"4C";
        when x"0FD5" => data_out<= x"8C";
        when x"0FD6" => data_out<= x"91";
        when x"0FD7" => data_out<= x"C9";
        when x"0FD8" => data_out<= x"BA";
        when x"0FD9" => data_out<= x"D0";
        when x"0FDA" => data_out<= x"03";
        when x"0FDB" => data_out<= x"4C";
        when x"0FDC" => data_out<= x"0E";
        when x"0FDD" => data_out<= x"91";
        when x"0FDE" => data_out<= x"C9";
        when x"0FDF" => data_out<= x"C0";
        when x"0FE0" => data_out<= x"D0";
        when x"0FE1" => data_out<= x"03";
        when x"0FE2" => data_out<= x"4C";
        when x"0FE3" => data_out<= x"4D";
        when x"0FE4" => data_out<= x"91";
        when x"0FE5" => data_out<= x"C9";
        when x"0FE6" => data_out<= x"C8";
        when x"0FE7" => data_out<= x"D0";
        when x"0FE8" => data_out<= x"03";
        when x"0FE9" => data_out<= x"4C";
        when x"0FEA" => data_out<= x"A5";
        when x"0FEB" => data_out<= x"90";
        when x"0FEC" => data_out<= x"C9";
        when x"0FED" => data_out<= x"C9";
        when x"0FEE" => data_out<= x"D0";
        when x"0FEF" => data_out<= x"03";
        when x"0FF0" => data_out<= x"4C";
        when x"0FF1" => data_out<= x"3F";
        when x"0FF2" => data_out<= x"91";
        when x"0FF3" => data_out<= x"C9";
        when x"0FF4" => data_out<= x"CA";
        when x"0FF5" => data_out<= x"D0";
        when x"0FF6" => data_out<= x"03";
        when x"0FF7" => data_out<= x"4C";
        when x"0FF8" => data_out<= x"AC";
        when x"0FF9" => data_out<= x"90";
        when x"0FFA" => data_out<= x"C9";
        when x"0FFB" => data_out<= x"D0";
        when x"0FFC" => data_out<= x"D0";
        when x"0FFD" => data_out<= x"03";
        when x"0FFE" => data_out<= x"4C";
        when x"0FFF" => data_out<= x"69";
        when x"1000" => data_out<= x"91";
        when x"1001" => data_out<= x"C9";
        when x"1002" => data_out<= x"D8";
        when x"1003" => data_out<= x"D0";
        when x"1004" => data_out<= x"03";
        when x"1005" => data_out<= x"4C";
        when x"1006" => data_out<= x"C8";
        when x"1007" => data_out<= x"90";
        when x"1008" => data_out<= x"C9";
        when x"1009" => data_out<= x"E0";
        when x"100A" => data_out<= x"D0";
        when x"100B" => data_out<= x"03";
        when x"100C" => data_out<= x"4C";
        when x"100D" => data_out<= x"46";
        when x"100E" => data_out<= x"91";
        when x"100F" => data_out<= x"C9";
        when x"1010" => data_out<= x"E8";
        when x"1011" => data_out<= x"D0";
        when x"1012" => data_out<= x"03";
        when x"1013" => data_out<= x"4C";
        when x"1014" => data_out<= x"9E";
        when x"1015" => data_out<= x"90";
        when x"1016" => data_out<= x"C9";
        when x"1017" => data_out<= x"E9";
        when x"1018" => data_out<= x"D0";
        when x"1019" => data_out<= x"03";
        when x"101A" => data_out<= x"4C";
        when x"101B" => data_out<= x"38";
        when x"101C" => data_out<= x"91";
        when x"101D" => data_out<= x"C9";
        when x"101E" => data_out<= x"EA";
        when x"101F" => data_out<= x"D0";
        when x"1020" => data_out<= x"03";
        when x"1021" => data_out<= x"4C";
        when x"1022" => data_out<= x"E4";
        when x"1023" => data_out<= x"90";
        when x"1024" => data_out<= x"C9";
        when x"1025" => data_out<= x"F0";
        when x"1026" => data_out<= x"D0";
        when x"1027" => data_out<= x"03";
        when x"1028" => data_out<= x"4C";
        when x"1029" => data_out<= x"70";
        when x"102A" => data_out<= x"91";
        when x"102B" => data_out<= x"C9";
        when x"102C" => data_out<= x"F8";
        when x"102D" => data_out<= x"D0";
        when x"102E" => data_out<= x"03";
        when x"102F" => data_out<= x"4C";
        when x"1030" => data_out<= x"CF";
        when x"1031" => data_out<= x"90";
        when x"1032" => data_out<= x"4C";
        when x"1033" => data_out<= x"A1";
        when x"1034" => data_out<= x"91";
        when x"1035" => data_out<= x"A9";
        when x"1036" => data_out<= x"29";
        when x"1037" => data_out<= x"A2";
        when x"1038" => data_out<= x"BD";
        when x"1039" => data_out<= x"4C";
        when x"103A" => data_out<= x"05";
        when x"103B" => data_out<= x"AF";
        when x"103C" => data_out<= x"A9";
        when x"103D" => data_out<= x"25";
        when x"103E" => data_out<= x"A2";
        when x"103F" => data_out<= x"BD";
        when x"1040" => data_out<= x"4C";
        when x"1041" => data_out<= x"05";
        when x"1042" => data_out<= x"AF";
        when x"1043" => data_out<= x"A9";
        when x"1044" => data_out<= x"21";
        when x"1045" => data_out<= x"A2";
        when x"1046" => data_out<= x"BD";
        when x"1047" => data_out<= x"4C";
        when x"1048" => data_out<= x"05";
        when x"1049" => data_out<= x"AF";
        when x"104A" => data_out<= x"A9";
        when x"104B" => data_out<= x"1D";
        when x"104C" => data_out<= x"A2";
        when x"104D" => data_out<= x"BD";
        when x"104E" => data_out<= x"4C";
        when x"104F" => data_out<= x"05";
        when x"1050" => data_out<= x"AF";
        when x"1051" => data_out<= x"A9";
        when x"1052" => data_out<= x"19";
        when x"1053" => data_out<= x"A2";
        when x"1054" => data_out<= x"BD";
        when x"1055" => data_out<= x"4C";
        when x"1056" => data_out<= x"05";
        when x"1057" => data_out<= x"AF";
        when x"1058" => data_out<= x"A9";
        when x"1059" => data_out<= x"67";
        when x"105A" => data_out<= x"A2";
        when x"105B" => data_out<= x"BC";
        when x"105C" => data_out<= x"4C";
        when x"105D" => data_out<= x"05";
        when x"105E" => data_out<= x"AF";
        when x"105F" => data_out<= x"A9";
        when x"1060" => data_out<= x"90";
        when x"1061" => data_out<= x"A2";
        when x"1062" => data_out<= x"BC";
        when x"1063" => data_out<= x"4C";
        when x"1064" => data_out<= x"05";
        when x"1065" => data_out<= x"AF";
        when x"1066" => data_out<= x"A9";
        when x"1067" => data_out<= x"4F";
        when x"1068" => data_out<= x"A2";
        when x"1069" => data_out<= x"BC";
        when x"106A" => data_out<= x"4C";
        when x"106B" => data_out<= x"05";
        when x"106C" => data_out<= x"AF";
        when x"106D" => data_out<= x"A9";
        when x"106E" => data_out<= x"5B";
        when x"106F" => data_out<= x"A2";
        when x"1070" => data_out<= x"BC";
        when x"1071" => data_out<= x"4C";
        when x"1072" => data_out<= x"05";
        when x"1073" => data_out<= x"AF";
        when x"1074" => data_out<= x"A9";
        when x"1075" => data_out<= x"BD";
        when x"1076" => data_out<= x"A2";
        when x"1077" => data_out<= x"BC";
        when x"1078" => data_out<= x"4C";
        when x"1079" => data_out<= x"05";
        when x"107A" => data_out<= x"AF";
        when x"107B" => data_out<= x"A9";
        when x"107C" => data_out<= x"C2";
        when x"107D" => data_out<= x"A2";
        when x"107E" => data_out<= x"BC";
        when x"107F" => data_out<= x"4C";
        when x"1080" => data_out<= x"05";
        when x"1081" => data_out<= x"AF";
        when x"1082" => data_out<= x"A9";
        when x"1083" => data_out<= x"6D";
        when x"1084" => data_out<= x"A2";
        when x"1085" => data_out<= x"BC";
        when x"1086" => data_out<= x"4C";
        when x"1087" => data_out<= x"05";
        when x"1088" => data_out<= x"AF";
        when x"1089" => data_out<= x"A9";
        when x"108A" => data_out<= x"73";
        when x"108B" => data_out<= x"A2";
        when x"108C" => data_out<= x"BC";
        when x"108D" => data_out<= x"4C";
        when x"108E" => data_out<= x"05";
        when x"108F" => data_out<= x"AF";
        when x"1090" => data_out<= x"A9";
        when x"1091" => data_out<= x"79";
        when x"1092" => data_out<= x"A2";
        when x"1093" => data_out<= x"BC";
        when x"1094" => data_out<= x"4C";
        when x"1095" => data_out<= x"05";
        when x"1096" => data_out<= x"AF";
        when x"1097" => data_out<= x"A9";
        when x"1098" => data_out<= x"85";
        when x"1099" => data_out<= x"A2";
        when x"109A" => data_out<= x"BC";
        when x"109B" => data_out<= x"4C";
        when x"109C" => data_out<= x"05";
        when x"109D" => data_out<= x"AF";
        when x"109E" => data_out<= x"A9";
        when x"109F" => data_out<= x"E9";
        when x"10A0" => data_out<= x"A2";
        when x"10A1" => data_out<= x"BC";
        when x"10A2" => data_out<= x"4C";
        when x"10A3" => data_out<= x"05";
        when x"10A4" => data_out<= x"AF";
        when x"10A5" => data_out<= x"A9";
        when x"10A6" => data_out<= x"E5";
        when x"10A7" => data_out<= x"A2";
        when x"10A8" => data_out<= x"BC";
        when x"10A9" => data_out<= x"4C";
        when x"10AA" => data_out<= x"05";
        when x"10AB" => data_out<= x"AF";
        when x"10AC" => data_out<= x"A9";
        when x"10AD" => data_out<= x"79";
        when x"10AE" => data_out<= x"A2";
        when x"10AF" => data_out<= x"BD";
        when x"10B0" => data_out<= x"4C";
        when x"10B1" => data_out<= x"05";
        when x"10B2" => data_out<= x"AF";
        when x"10B3" => data_out<= x"A9";
        when x"10B4" => data_out<= x"ED";
        when x"10B5" => data_out<= x"A2";
        when x"10B6" => data_out<= x"BC";
        when x"10B7" => data_out<= x"4C";
        when x"10B8" => data_out<= x"05";
        when x"10B9" => data_out<= x"AF";
        when x"10BA" => data_out<= x"A9";
        when x"10BB" => data_out<= x"F1";
        when x"10BC" => data_out<= x"A2";
        when x"10BD" => data_out<= x"BC";
        when x"10BE" => data_out<= x"4C";
        when x"10BF" => data_out<= x"05";
        when x"10C0" => data_out<= x"AF";
        when x"10C1" => data_out<= x"A9";
        when x"10C2" => data_out<= x"F5";
        when x"10C3" => data_out<= x"A2";
        when x"10C4" => data_out<= x"BC";
        when x"10C5" => data_out<= x"4C";
        when x"10C6" => data_out<= x"05";
        when x"10C7" => data_out<= x"AF";
        when x"10C8" => data_out<= x"A9";
        when x"10C9" => data_out<= x"F9";
        when x"10CA" => data_out<= x"A2";
        when x"10CB" => data_out<= x"BC";
        when x"10CC" => data_out<= x"4C";
        when x"10CD" => data_out<= x"05";
        when x"10CE" => data_out<= x"AF";
        when x"10CF" => data_out<= x"A9";
        when x"10D0" => data_out<= x"FD";
        when x"10D1" => data_out<= x"A2";
        when x"10D2" => data_out<= x"BC";
        when x"10D3" => data_out<= x"4C";
        when x"10D4" => data_out<= x"05";
        when x"10D5" => data_out<= x"AF";
        when x"10D6" => data_out<= x"A9";
        when x"10D7" => data_out<= x"15";
        when x"10D8" => data_out<= x"A2";
        when x"10D9" => data_out<= x"BD";
        when x"10DA" => data_out<= x"4C";
        when x"10DB" => data_out<= x"05";
        when x"10DC" => data_out<= x"AF";
        when x"10DD" => data_out<= x"A9";
        when x"10DE" => data_out<= x"35";
        when x"10DF" => data_out<= x"A2";
        when x"10E0" => data_out<= x"BD";
        when x"10E1" => data_out<= x"4C";
        when x"10E2" => data_out<= x"05";
        when x"10E3" => data_out<= x"AF";
        when x"10E4" => data_out<= x"A9";
        when x"10E5" => data_out<= x"3D";
        when x"10E6" => data_out<= x"A2";
        when x"10E7" => data_out<= x"BD";
        when x"10E8" => data_out<= x"4C";
        when x"10E9" => data_out<= x"05";
        when x"10EA" => data_out<= x"AF";
        when x"10EB" => data_out<= x"A9";
        when x"10EC" => data_out<= x"41";
        when x"10ED" => data_out<= x"A2";
        when x"10EE" => data_out<= x"BD";
        when x"10EF" => data_out<= x"4C";
        when x"10F0" => data_out<= x"05";
        when x"10F1" => data_out<= x"AF";
        when x"10F2" => data_out<= x"A9";
        when x"10F3" => data_out<= x"49";
        when x"10F4" => data_out<= x"A2";
        when x"10F5" => data_out<= x"BD";
        when x"10F6" => data_out<= x"4C";
        when x"10F7" => data_out<= x"05";
        when x"10F8" => data_out<= x"AF";
        when x"10F9" => data_out<= x"A9";
        when x"10FA" => data_out<= x"4D";
        when x"10FB" => data_out<= x"A2";
        when x"10FC" => data_out<= x"BD";
        when x"10FD" => data_out<= x"4C";
        when x"10FE" => data_out<= x"05";
        when x"10FF" => data_out<= x"AF";
        when x"1100" => data_out<= x"A9";
        when x"1101" => data_out<= x"51";
        when x"1102" => data_out<= x"A2";
        when x"1103" => data_out<= x"BD";
        when x"1104" => data_out<= x"4C";
        when x"1105" => data_out<= x"05";
        when x"1106" => data_out<= x"AF";
        when x"1107" => data_out<= x"A9";
        when x"1108" => data_out<= x"5D";
        when x"1109" => data_out<= x"A2";
        when x"110A" => data_out<= x"BD";
        when x"110B" => data_out<= x"4C";
        when x"110C" => data_out<= x"05";
        when x"110D" => data_out<= x"AF";
        when x"110E" => data_out<= x"A9";
        when x"110F" => data_out<= x"65";
        when x"1110" => data_out<= x"A2";
        when x"1111" => data_out<= x"BD";
        when x"1112" => data_out<= x"4C";
        when x"1113" => data_out<= x"05";
        when x"1114" => data_out<= x"AF";
        when x"1115" => data_out<= x"A9";
        when x"1116" => data_out<= x"69";
        when x"1117" => data_out<= x"A2";
        when x"1118" => data_out<= x"BD";
        when x"1119" => data_out<= x"4C";
        when x"111A" => data_out<= x"05";
        when x"111B" => data_out<= x"AF";
        when x"111C" => data_out<= x"A9";
        when x"111D" => data_out<= x"6D";
        when x"111E" => data_out<= x"A2";
        when x"111F" => data_out<= x"BD";
        when x"1120" => data_out<= x"4C";
        when x"1121" => data_out<= x"05";
        when x"1122" => data_out<= x"AF";
        when x"1123" => data_out<= x"A9";
        when x"1124" => data_out<= x"71";
        when x"1125" => data_out<= x"A2";
        when x"1126" => data_out<= x"BD";
        when x"1127" => data_out<= x"4C";
        when x"1128" => data_out<= x"05";
        when x"1129" => data_out<= x"AF";
        when x"112A" => data_out<= x"A9";
        when x"112B" => data_out<= x"75";
        when x"112C" => data_out<= x"A2";
        when x"112D" => data_out<= x"BD";
        when x"112E" => data_out<= x"4C";
        when x"112F" => data_out<= x"05";
        when x"1130" => data_out<= x"AF";
        when x"1131" => data_out<= x"A9";
        when x"1132" => data_out<= x"A9";
        when x"1133" => data_out<= x"A2";
        when x"1134" => data_out<= x"BC";
        when x"1135" => data_out<= x"4C";
        when x"1136" => data_out<= x"05";
        when x"1137" => data_out<= x"AF";
        when x"1138" => data_out<= x"A9";
        when x"1139" => data_out<= x"E0";
        when x"113A" => data_out<= x"A2";
        when x"113B" => data_out<= x"BC";
        when x"113C" => data_out<= x"4C";
        when x"113D" => data_out<= x"05";
        when x"113E" => data_out<= x"AF";
        when x"113F" => data_out<= x"A9";
        when x"1140" => data_out<= x"DB";
        when x"1141" => data_out<= x"A2";
        when x"1142" => data_out<= x"BC";
        when x"1143" => data_out<= x"4C";
        when x"1144" => data_out<= x"05";
        when x"1145" => data_out<= x"AF";
        when x"1146" => data_out<= x"A9";
        when x"1147" => data_out<= x"D6";
        when x"1148" => data_out<= x"A2";
        when x"1149" => data_out<= x"BC";
        when x"114A" => data_out<= x"4C";
        when x"114B" => data_out<= x"05";
        when x"114C" => data_out<= x"AF";
        when x"114D" => data_out<= x"A9";
        when x"114E" => data_out<= x"D1";
        when x"114F" => data_out<= x"A2";
        when x"1150" => data_out<= x"BC";
        when x"1151" => data_out<= x"4C";
        when x"1152" => data_out<= x"05";
        when x"1153" => data_out<= x"AF";
        when x"1154" => data_out<= x"A9";
        when x"1155" => data_out<= x"CC";
        when x"1156" => data_out<= x"A2";
        when x"1157" => data_out<= x"BC";
        when x"1158" => data_out<= x"4C";
        when x"1159" => data_out<= x"05";
        when x"115A" => data_out<= x"AF";
        when x"115B" => data_out<= x"A9";
        when x"115C" => data_out<= x"B3";
        when x"115D" => data_out<= x"A2";
        when x"115E" => data_out<= x"BC";
        when x"115F" => data_out<= x"4C";
        when x"1160" => data_out<= x"05";
        when x"1161" => data_out<= x"AF";
        when x"1162" => data_out<= x"A9";
        when x"1163" => data_out<= x"AE";
        when x"1164" => data_out<= x"A2";
        when x"1165" => data_out<= x"BC";
        when x"1166" => data_out<= x"4C";
        when x"1167" => data_out<= x"05";
        when x"1168" => data_out<= x"AF";
        when x"1169" => data_out<= x"A9";
        when x"116A" => data_out<= x"05";
        when x"116B" => data_out<= x"A2";
        when x"116C" => data_out<= x"BD";
        when x"116D" => data_out<= x"4C";
        when x"116E" => data_out<= x"05";
        when x"116F" => data_out<= x"AF";
        when x"1170" => data_out<= x"A9";
        when x"1171" => data_out<= x"09";
        when x"1172" => data_out<= x"A2";
        when x"1173" => data_out<= x"BD";
        when x"1174" => data_out<= x"4C";
        when x"1175" => data_out<= x"05";
        when x"1176" => data_out<= x"AF";
        when x"1177" => data_out<= x"A9";
        when x"1178" => data_out<= x"0D";
        when x"1179" => data_out<= x"A2";
        when x"117A" => data_out<= x"BD";
        when x"117B" => data_out<= x"4C";
        when x"117C" => data_out<= x"05";
        when x"117D" => data_out<= x"AF";
        when x"117E" => data_out<= x"A9";
        when x"117F" => data_out<= x"2D";
        when x"1180" => data_out<= x"A2";
        when x"1181" => data_out<= x"BD";
        when x"1182" => data_out<= x"4C";
        when x"1183" => data_out<= x"05";
        when x"1184" => data_out<= x"AF";
        when x"1185" => data_out<= x"A9";
        when x"1186" => data_out<= x"31";
        when x"1187" => data_out<= x"A2";
        when x"1188" => data_out<= x"BD";
        when x"1189" => data_out<= x"4C";
        when x"118A" => data_out<= x"05";
        when x"118B" => data_out<= x"AF";
        when x"118C" => data_out<= x"A9";
        when x"118D" => data_out<= x"45";
        when x"118E" => data_out<= x"A2";
        when x"118F" => data_out<= x"BD";
        when x"1190" => data_out<= x"4C";
        when x"1191" => data_out<= x"05";
        when x"1192" => data_out<= x"AF";
        when x"1193" => data_out<= x"A9";
        when x"1194" => data_out<= x"55";
        when x"1195" => data_out<= x"A2";
        when x"1196" => data_out<= x"BD";
        when x"1197" => data_out<= x"4C";
        when x"1198" => data_out<= x"05";
        when x"1199" => data_out<= x"AF";
        when x"119A" => data_out<= x"A9";
        when x"119B" => data_out<= x"59";
        when x"119C" => data_out<= x"A2";
        when x"119D" => data_out<= x"BD";
        when x"119E" => data_out<= x"4C";
        when x"119F" => data_out<= x"05";
        when x"11A0" => data_out<= x"AF";
        when x"11A1" => data_out<= x"A9";
        when x"11A2" => data_out<= x"61";
        when x"11A3" => data_out<= x"A2";
        when x"11A4" => data_out<= x"BD";
        when x"11A5" => data_out<= x"4C";
        when x"11A6" => data_out<= x"05";
        when x"11A7" => data_out<= x"AF";
        when x"11A8" => data_out<= x"20";
        when x"11A9" => data_out<= x"65";
        when x"11AA" => data_out<= x"B0";
        when x"11AB" => data_out<= x"A0";
        when x"11AC" => data_out<= x"00";
        when x"11AD" => data_out<= x"B1";
        when x"11AE" => data_out<= x"0C";
        when x"11AF" => data_out<= x"F0";
        when x"11B0" => data_out<= x"5C";
        when x"11B1" => data_out<= x"C9";
        when x"11B2" => data_out<= x"40";
        when x"11B3" => data_out<= x"F0";
        when x"11B4" => data_out<= x"58";
        when x"11B5" => data_out<= x"C9";
        when x"11B6" => data_out<= x"60";
        when x"11B7" => data_out<= x"F0";
        when x"11B8" => data_out<= x"54";
        when x"11B9" => data_out<= x"C9";
        when x"11BA" => data_out<= x"E8";
        when x"11BB" => data_out<= x"F0";
        when x"11BC" => data_out<= x"50";
        when x"11BD" => data_out<= x"C9";
        when x"11BE" => data_out<= x"C8";
        when x"11BF" => data_out<= x"F0";
        when x"11C0" => data_out<= x"4C";
        when x"11C1" => data_out<= x"C9";
        when x"11C2" => data_out<= x"CA";
        when x"11C3" => data_out<= x"F0";
        when x"11C4" => data_out<= x"48";
        when x"11C5" => data_out<= x"C9";
        when x"11C6" => data_out<= x"88";
        when x"11C7" => data_out<= x"F0";
        when x"11C8" => data_out<= x"44";
        when x"11C9" => data_out<= x"C9";
        when x"11CA" => data_out<= x"18";
        when x"11CB" => data_out<= x"F0";
        when x"11CC" => data_out<= x"40";
        when x"11CD" => data_out<= x"C9";
        when x"11CE" => data_out<= x"38";
        when x"11CF" => data_out<= x"F0";
        when x"11D0" => data_out<= x"3C";
        when x"11D1" => data_out<= x"C9";
        when x"11D2" => data_out<= x"D8";
        when x"11D3" => data_out<= x"F0";
        when x"11D4" => data_out<= x"38";
        when x"11D5" => data_out<= x"C9";
        when x"11D6" => data_out<= x"F8";
        when x"11D7" => data_out<= x"F0";
        when x"11D8" => data_out<= x"34";
        when x"11D9" => data_out<= x"C9";
        when x"11DA" => data_out<= x"58";
        when x"11DB" => data_out<= x"F0";
        when x"11DC" => data_out<= x"30";
        when x"11DD" => data_out<= x"C9";
        when x"11DE" => data_out<= x"78";
        when x"11DF" => data_out<= x"F0";
        when x"11E0" => data_out<= x"2C";
        when x"11E1" => data_out<= x"C9";
        when x"11E2" => data_out<= x"EA";
        when x"11E3" => data_out<= x"F0";
        when x"11E4" => data_out<= x"28";
        when x"11E5" => data_out<= x"C9";
        when x"11E6" => data_out<= x"AA";
        when x"11E7" => data_out<= x"F0";
        when x"11E8" => data_out<= x"24";
        when x"11E9" => data_out<= x"C9";
        when x"11EA" => data_out<= x"A8";
        when x"11EB" => data_out<= x"F0";
        when x"11EC" => data_out<= x"20";
        when x"11ED" => data_out<= x"C9";
        when x"11EE" => data_out<= x"8A";
        when x"11EF" => data_out<= x"F0";
        when x"11F0" => data_out<= x"1C";
        when x"11F1" => data_out<= x"C9";
        when x"11F2" => data_out<= x"98";
        when x"11F3" => data_out<= x"F0";
        when x"11F4" => data_out<= x"18";
        when x"11F5" => data_out<= x"C9";
        when x"11F6" => data_out<= x"9A";
        when x"11F7" => data_out<= x"F0";
        when x"11F8" => data_out<= x"14";
        when x"11F9" => data_out<= x"C9";
        when x"11FA" => data_out<= x"BA";
        when x"11FB" => data_out<= x"F0";
        when x"11FC" => data_out<= x"10";
        when x"11FD" => data_out<= x"C9";
        when x"11FE" => data_out<= x"48";
        when x"11FF" => data_out<= x"F0";
        when x"1200" => data_out<= x"0C";
        when x"1201" => data_out<= x"C9";
        when x"1202" => data_out<= x"68";
        when x"1203" => data_out<= x"F0";
        when x"1204" => data_out<= x"08";
        when x"1205" => data_out<= x"C9";
        when x"1206" => data_out<= x"08";
        when x"1207" => data_out<= x"F0";
        when x"1208" => data_out<= x"04";
        when x"1209" => data_out<= x"C9";
        when x"120A" => data_out<= x"28";
        when x"120B" => data_out<= x"D0";
        when x"120C" => data_out<= x"07";
        when x"120D" => data_out<= x"A2";
        when x"120E" => data_out<= x"00";
        when x"120F" => data_out<= x"A9";
        when x"1210" => data_out<= x"01";
        when x"1211" => data_out<= x"4C";
        when x"1212" => data_out<= x"05";
        when x"1213" => data_out<= x"AF";
        when x"1214" => data_out<= x"B1";
        when x"1215" => data_out<= x"0C";
        when x"1216" => data_out<= x"29";
        when x"1217" => data_out<= x"0F";
        when x"1218" => data_out<= x"C9";
        when x"1219" => data_out<= x"09";
        when x"121A" => data_out<= x"F0";
        when x"121B" => data_out<= x"2A";
        when x"121C" => data_out<= x"B1";
        when x"121D" => data_out<= x"0C";
        when x"121E" => data_out<= x"29";
        when x"121F" => data_out<= x"0F";
        when x"1220" => data_out<= x"C9";
        when x"1221" => data_out<= x"05";
        when x"1222" => data_out<= x"F0";
        when x"1223" => data_out<= x"22";
        when x"1224" => data_out<= x"B1";
        when x"1225" => data_out<= x"0C";
        when x"1226" => data_out<= x"29";
        when x"1227" => data_out<= x"0F";
        when x"1228" => data_out<= x"C9";
        when x"1229" => data_out<= x"06";
        when x"122A" => data_out<= x"F0";
        when x"122B" => data_out<= x"1A";
        when x"122C" => data_out<= x"B1";
        when x"122D" => data_out<= x"0C";
        when x"122E" => data_out<= x"29";
        when x"122F" => data_out<= x"1F";
        when x"1230" => data_out<= x"C9";
        when x"1231" => data_out<= x"10";
        when x"1232" => data_out<= x"F0";
        when x"1233" => data_out<= x"12";
        when x"1234" => data_out<= x"B1";
        when x"1235" => data_out<= x"0C";
        when x"1236" => data_out<= x"C9";
        when x"1237" => data_out<= x"A2";
        when x"1238" => data_out<= x"F0";
        when x"1239" => data_out<= x"0C";
        when x"123A" => data_out<= x"C9";
        when x"123B" => data_out<= x"A0";
        when x"123C" => data_out<= x"F0";
        when x"123D" => data_out<= x"08";
        when x"123E" => data_out<= x"C9";
        when x"123F" => data_out<= x"E0";
        when x"1240" => data_out<= x"F0";
        when x"1241" => data_out<= x"04";
        when x"1242" => data_out<= x"C9";
        when x"1243" => data_out<= x"C0";
        when x"1244" => data_out<= x"D0";
        when x"1245" => data_out<= x"05";
        when x"1246" => data_out<= x"A2";
        when x"1247" => data_out<= x"00";
        when x"1248" => data_out<= x"4C";
        when x"1249" => data_out<= x"73";
        when x"124A" => data_out<= x"92";
        when x"124B" => data_out<= x"B1";
        when x"124C" => data_out<= x"0C";
        when x"124D" => data_out<= x"C9";
        when x"124E" => data_out<= x"20";
        when x"124F" => data_out<= x"F0";
        when x"1250" => data_out<= x"1B";
        when x"1251" => data_out<= x"C9";
        when x"1252" => data_out<= x"4C";
        when x"1253" => data_out<= x"F0";
        when x"1254" => data_out<= x"17";
        when x"1255" => data_out<= x"C9";
        when x"1256" => data_out<= x"6C";
        when x"1257" => data_out<= x"F0";
        when x"1258" => data_out<= x"13";
        when x"1259" => data_out<= x"29";
        when x"125A" => data_out<= x"0F";
        when x"125B" => data_out<= x"C9";
        when x"125C" => data_out<= x"0D";
        when x"125D" => data_out<= x"F0";
        when x"125E" => data_out<= x"0D";
        when x"125F" => data_out<= x"B1";
        when x"1260" => data_out<= x"0C";
        when x"1261" => data_out<= x"29";
        when x"1262" => data_out<= x"0F";
        when x"1263" => data_out<= x"C9";
        when x"1264" => data_out<= x"0E";
        when x"1265" => data_out<= x"F0";
        when x"1266" => data_out<= x"05";
        when x"1267" => data_out<= x"A2";
        when x"1268" => data_out<= x"00";
        when x"1269" => data_out<= x"4C";
        when x"126A" => data_out<= x"73";
        when x"126B" => data_out<= x"92";
        when x"126C" => data_out<= x"A2";
        when x"126D" => data_out<= x"00";
        when x"126E" => data_out<= x"A9";
        when x"126F" => data_out<= x"03";
        when x"1270" => data_out<= x"4C";
        when x"1271" => data_out<= x"05";
        when x"1272" => data_out<= x"AF";
        when x"1273" => data_out<= x"A9";
        when x"1274" => data_out<= x"02";
        when x"1275" => data_out<= x"4C";
        when x"1276" => data_out<= x"05";
        when x"1277" => data_out<= x"AF";
        when x"1278" => data_out<= x"20";
        when x"1279" => data_out<= x"65";
        when x"127A" => data_out<= x"B0";
        when x"127B" => data_out<= x"20";
        when x"127C" => data_out<= x"A7";
        when x"127D" => data_out<= x"AE";
        when x"127E" => data_out<= x"A9";
        when x"127F" => data_out<= x"00";
        when x"1280" => data_out<= x"A0";
        when x"1281" => data_out<= x"06";
        when x"1282" => data_out<= x"91";
        when x"1283" => data_out<= x"0C";
        when x"1284" => data_out<= x"C8";
        when x"1285" => data_out<= x"D1";
        when x"1286" => data_out<= x"0C";
        when x"1287" => data_out<= x"90";
        when x"1288" => data_out<= x"03";
        when x"1289" => data_out<= x"4C";
        when x"128A" => data_out<= x"76";
        when x"128B" => data_out<= x"93";
        when x"128C" => data_out<= x"A0";
        when x"128D" => data_out<= x"09";
        when x"128E" => data_out<= x"20";
        when x"128F" => data_out<= x"4F";
        when x"1290" => data_out<= x"AF";
        when x"1291" => data_out<= x"20";
        when x"1292" => data_out<= x"49";
        when x"1293" => data_out<= x"89";
        when x"1294" => data_out<= x"A0";
        when x"1295" => data_out<= x"03";
        when x"1296" => data_out<= x"91";
        when x"1297" => data_out<= x"0C";
        when x"1298" => data_out<= x"20";
        when x"1299" => data_out<= x"A8";
        when x"129A" => data_out<= x"91";
        when x"129B" => data_out<= x"A0";
        when x"129C" => data_out<= x"04";
        when x"129D" => data_out<= x"91";
        when x"129E" => data_out<= x"0C";
        when x"129F" => data_out<= x"A9";
        when x"12A0" => data_out<= x"00";
        when x"12A1" => data_out<= x"C8";
        when x"12A2" => data_out<= x"91";
        when x"12A3" => data_out<= x"0C";
        when x"12A4" => data_out<= x"88";
        when x"12A5" => data_out<= x"D1";
        when x"12A6" => data_out<= x"0C";
        when x"12A7" => data_out<= x"B0";
        when x"12A8" => data_out<= x"31";
        when x"12A9" => data_out<= x"A5";
        when x"12AA" => data_out<= x"0C";
        when x"12AB" => data_out<= x"A6";
        when x"12AC" => data_out<= x"0D";
        when x"12AD" => data_out<= x"C8";
        when x"12AE" => data_out<= x"18";
        when x"12AF" => data_out<= x"71";
        when x"12B0" => data_out<= x"0C";
        when x"12B1" => data_out<= x"90";
        when x"12B2" => data_out<= x"01";
        when x"12B3" => data_out<= x"E8";
        when x"12B4" => data_out<= x"20";
        when x"12B5" => data_out<= x"7B";
        when x"12B6" => data_out<= x"B0";
        when x"12B7" => data_out<= x"A0";
        when x"12B8" => data_out<= x"07";
        when x"12B9" => data_out<= x"B1";
        when x"12BA" => data_out<= x"0C";
        when x"12BB" => data_out<= x"18";
        when x"12BC" => data_out<= x"A0";
        when x"12BD" => data_out<= x"0A";
        when x"12BE" => data_out<= x"71";
        when x"12BF" => data_out<= x"0C";
        when x"12C0" => data_out<= x"48";
        when x"12C1" => data_out<= x"A9";
        when x"12C2" => data_out<= x"00";
        when x"12C3" => data_out<= x"C8";
        when x"12C4" => data_out<= x"71";
        when x"12C5" => data_out<= x"0C";
        when x"12C6" => data_out<= x"AA";
        when x"12C7" => data_out<= x"68";
        when x"12C8" => data_out<= x"20";
        when x"12C9" => data_out<= x"49";
        when x"12CA" => data_out<= x"89";
        when x"12CB" => data_out<= x"A0";
        when x"12CC" => data_out<= x"00";
        when x"12CD" => data_out<= x"20";
        when x"12CE" => data_out<= x"AD";
        when x"12CF" => data_out<= x"B0";
        when x"12D0" => data_out<= x"A0";
        when x"12D1" => data_out<= x"05";
        when x"12D2" => data_out<= x"B1";
        when x"12D3" => data_out<= x"0C";
        when x"12D4" => data_out<= x"18";
        when x"12D5" => data_out<= x"69";
        when x"12D6" => data_out<= x"01";
        when x"12D7" => data_out<= x"4C";
        when x"12D8" => data_out<= x"A2";
        when x"12D9" => data_out<= x"92";
        when x"12DA" => data_out<= x"A0";
        when x"12DB" => data_out<= x"09";
        when x"12DC" => data_out<= x"20";
        when x"12DD" => data_out<= x"4F";
        when x"12DE" => data_out<= x"AF";
        when x"12DF" => data_out<= x"20";
        when x"12E0" => data_out<= x"31";
        when x"12E1" => data_out<= x"8C";
        when x"12E2" => data_out<= x"A9";
        when x"12E3" => data_out<= x"02";
        when x"12E4" => data_out<= x"A2";
        when x"12E5" => data_out<= x"BD";
        when x"12E6" => data_out<= x"20";
        when x"12E7" => data_out<= x"22";
        when x"12E8" => data_out<= x"81";
        when x"12E9" => data_out<= x"A9";
        when x"12EA" => data_out<= x"00";
        when x"12EB" => data_out<= x"A0";
        when x"12EC" => data_out<= x"05";
        when x"12ED" => data_out<= x"91";
        when x"12EE" => data_out<= x"0C";
        when x"12EF" => data_out<= x"C9";
        when x"12F0" => data_out<= x"03";
        when x"12F1" => data_out<= x"B0";
        when x"12F2" => data_out<= x"34";
        when x"12F3" => data_out<= x"B1";
        when x"12F4" => data_out<= x"0C";
        when x"12F5" => data_out<= x"88";
        when x"12F6" => data_out<= x"D1";
        when x"12F7" => data_out<= x"0C";
        when x"12F8" => data_out<= x"B0";
        when x"12F9" => data_out<= x"19";
        when x"12FA" => data_out<= x"A5";
        when x"12FB" => data_out<= x"0C";
        when x"12FC" => data_out<= x"A6";
        when x"12FD" => data_out<= x"0D";
        when x"12FE" => data_out<= x"C8";
        when x"12FF" => data_out<= x"18";
        when x"1300" => data_out<= x"71";
        when x"1301" => data_out<= x"0C";
        when x"1302" => data_out<= x"90";
        when x"1303" => data_out<= x"01";
        when x"1304" => data_out<= x"E8";
        when x"1305" => data_out<= x"85";
        when x"1306" => data_out<= x"14";
        when x"1307" => data_out<= x"86";
        when x"1308" => data_out<= x"15";
        when x"1309" => data_out<= x"A0";
        when x"130A" => data_out<= x"00";
        when x"130B" => data_out<= x"B1";
        when x"130C" => data_out<= x"14";
        when x"130D" => data_out<= x"20";
        when x"130E" => data_out<= x"FD";
        when x"130F" => data_out<= x"8B";
        when x"1310" => data_out<= x"4C";
        when x"1311" => data_out<= x"1A";
        when x"1312" => data_out<= x"93";
        when x"1313" => data_out<= x"A9";
        when x"1314" => data_out<= x"02";
        when x"1315" => data_out<= x"A2";
        when x"1316" => data_out<= x"BD";
        when x"1317" => data_out<= x"20";
        when x"1318" => data_out<= x"22";
        when x"1319" => data_out<= x"81";
        when x"131A" => data_out<= x"20";
        when x"131B" => data_out<= x"8C";
        when x"131C" => data_out<= x"8C";
        when x"131D" => data_out<= x"A0";
        when x"131E" => data_out<= x"05";
        when x"131F" => data_out<= x"B1";
        when x"1320" => data_out<= x"0C";
        when x"1321" => data_out<= x"18";
        when x"1322" => data_out<= x"69";
        when x"1323" => data_out<= x"01";
        when x"1324" => data_out<= x"4C";
        when x"1325" => data_out<= x"ED";
        when x"1326" => data_out<= x"92";
        when x"1327" => data_out<= x"A0";
        when x"1328" => data_out<= x"03";
        when x"1329" => data_out<= x"B1";
        when x"132A" => data_out<= x"0C";
        when x"132B" => data_out<= x"20";
        when x"132C" => data_out<= x"C1";
        when x"132D" => data_out<= x"8E";
        when x"132E" => data_out<= x"20";
        when x"132F" => data_out<= x"22";
        when x"1330" => data_out<= x"81";
        when x"1331" => data_out<= x"A0";
        when x"1332" => data_out<= x"04";
        when x"1333" => data_out<= x"B1";
        when x"1334" => data_out<= x"0C";
        when x"1335" => data_out<= x"C9";
        when x"1336" => data_out<= x"02";
        when x"1337" => data_out<= x"D0";
        when x"1338" => data_out<= x"0A";
        when x"1339" => data_out<= x"A9";
        when x"133A" => data_out<= x"0F";
        when x"133B" => data_out<= x"A2";
        when x"133C" => data_out<= x"B9";
        when x"133D" => data_out<= x"20";
        when x"133E" => data_out<= x"22";
        when x"133F" => data_out<= x"81";
        when x"1340" => data_out<= x"4C";
        when x"1341" => data_out<= x"57";
        when x"1342" => data_out<= x"93";
        when x"1343" => data_out<= x"B1";
        when x"1344" => data_out<= x"0C";
        when x"1345" => data_out<= x"C9";
        when x"1346" => data_out<= x"03";
        when x"1347" => data_out<= x"D0";
        when x"1348" => data_out<= x"15";
        when x"1349" => data_out<= x"A9";
        when x"134A" => data_out<= x"0F";
        when x"134B" => data_out<= x"A2";
        when x"134C" => data_out<= x"B9";
        when x"134D" => data_out<= x"20";
        when x"134E" => data_out<= x"22";
        when x"134F" => data_out<= x"81";
        when x"1350" => data_out<= x"A0";
        when x"1351" => data_out<= x"02";
        when x"1352" => data_out<= x"B1";
        when x"1353" => data_out<= x"0C";
        when x"1354" => data_out<= x"20";
        when x"1355" => data_out<= x"FD";
        when x"1356" => data_out<= x"8B";
        when x"1357" => data_out<= x"A0";
        when x"1358" => data_out<= x"01";
        when x"1359" => data_out<= x"B1";
        when x"135A" => data_out<= x"0C";
        when x"135B" => data_out<= x"20";
        when x"135C" => data_out<= x"FD";
        when x"135D" => data_out<= x"8B";
        when x"135E" => data_out<= x"20";
        when x"135F" => data_out<= x"45";
        when x"1360" => data_out<= x"8C";
        when x"1361" => data_out<= x"A0";
        when x"1362" => data_out<= x"04";
        when x"1363" => data_out<= x"B1";
        when x"1364" => data_out<= x"0C";
        when x"1365" => data_out<= x"A2";
        when x"1366" => data_out<= x"00";
        when x"1367" => data_out<= x"A0";
        when x"1368" => data_out<= x"08";
        when x"1369" => data_out<= x"20";
        when x"136A" => data_out<= x"04";
        when x"136B" => data_out<= x"AE";
        when x"136C" => data_out<= x"A0";
        when x"136D" => data_out<= x"06";
        when x"136E" => data_out<= x"B1";
        when x"136F" => data_out<= x"0C";
        when x"1370" => data_out<= x"18";
        when x"1371" => data_out<= x"69";
        when x"1372" => data_out<= x"01";
        when x"1373" => data_out<= x"4C";
        when x"1374" => data_out<= x"82";
        when x"1375" => data_out<= x"92";
        when x"1376" => data_out<= x"A0";
        when x"1377" => data_out<= x"09";
        when x"1378" => data_out<= x"20";
        when x"1379" => data_out<= x"4F";
        when x"137A" => data_out<= x"AF";
        when x"137B" => data_out<= x"8D";
        when x"137C" => data_out<= x"00";
        when x"137D" => data_out<= x"02";
        when x"137E" => data_out<= x"8E";
        when x"137F" => data_out<= x"01";
        when x"1380" => data_out<= x"02";
        when x"1381" => data_out<= x"A0";
        when x"1382" => data_out<= x"0A";
        when x"1383" => data_out<= x"4C";
        when x"1384" => data_out<= x"14";
        when x"1385" => data_out<= x"AE";
        when x"1386" => data_out<= x"20";
        when x"1387" => data_out<= x"7B";
        when x"1388" => data_out<= x"B0";
        when x"1389" => data_out<= x"20";
        when x"138A" => data_out<= x"9A";
        when x"138B" => data_out<= x"AE";
        when x"138C" => data_out<= x"A9";
        when x"138D" => data_out<= x"00";
        when x"138E" => data_out<= x"20";
        when x"138F" => data_out<= x"65";
        when x"1390" => data_out<= x"B0";
        when x"1391" => data_out<= x"A0";
        when x"1392" => data_out<= x"07";
        when x"1393" => data_out<= x"B1";
        when x"1394" => data_out<= x"0C";
        when x"1395" => data_out<= x"C8";
        when x"1396" => data_out<= x"11";
        when x"1397" => data_out<= x"0C";
        when x"1398" => data_out<= x"D0";
        when x"1399" => data_out<= x"4A";
        when x"139A" => data_out<= x"A9";
        when x"139B" => data_out<= x"30";
        when x"139C" => data_out<= x"20";
        when x"139D" => data_out<= x"F0";
        when x"139E" => data_out<= x"80";
        when x"139F" => data_out<= x"4C";
        when x"13A0" => data_out<= x"17";
        when x"13A1" => data_out<= x"94";
        when x"13A2" => data_out<= x"A0";
        when x"13A3" => data_out<= x"00";
        when x"13A4" => data_out<= x"A2";
        when x"13A5" => data_out<= x"00";
        when x"13A6" => data_out<= x"B1";
        when x"13A7" => data_out<= x"0C";
        when x"13A8" => data_out<= x"48";
        when x"13A9" => data_out<= x"18";
        when x"13AA" => data_out<= x"69";
        when x"13AB" => data_out<= x"01";
        when x"13AC" => data_out<= x"91";
        when x"13AD" => data_out<= x"0C";
        when x"13AE" => data_out<= x"68";
        when x"13AF" => data_out<= x"18";
        when x"13B0" => data_out<= x"69";
        when x"13B1" => data_out<= x"01";
        when x"13B2" => data_out<= x"90";
        when x"13B3" => data_out<= x"02";
        when x"13B4" => data_out<= x"E8";
        when x"13B5" => data_out<= x"18";
        when x"13B6" => data_out<= x"65";
        when x"13B7" => data_out<= x"0C";
        when x"13B8" => data_out<= x"A8";
        when x"13B9" => data_out<= x"8A";
        when x"13BA" => data_out<= x"65";
        when x"13BB" => data_out<= x"0D";
        when x"13BC" => data_out<= x"AA";
        when x"13BD" => data_out<= x"98";
        when x"13BE" => data_out<= x"20";
        when x"13BF" => data_out<= x"7B";
        when x"13C0" => data_out<= x"B0";
        when x"13C1" => data_out<= x"A0";
        when x"13C2" => data_out<= x"0C";
        when x"13C3" => data_out<= x"20";
        when x"13C4" => data_out<= x"93";
        when x"13C5" => data_out<= x"B0";
        when x"13C6" => data_out<= x"A9";
        when x"13C7" => data_out<= x"0A";
        when x"13C8" => data_out<= x"20";
        when x"13C9" => data_out<= x"6F";
        when x"13CA" => data_out<= x"B1";
        when x"13CB" => data_out<= x"A0";
        when x"13CC" => data_out<= x"30";
        when x"13CD" => data_out<= x"20";
        when x"13CE" => data_out<= x"FC";
        when x"13CF" => data_out<= x"AE";
        when x"13D0" => data_out<= x"A0";
        when x"13D1" => data_out<= x"00";
        when x"13D2" => data_out<= x"20";
        when x"13D3" => data_out<= x"AD";
        when x"13D4" => data_out<= x"B0";
        when x"13D5" => data_out<= x"A0";
        when x"13D6" => data_out<= x"0A";
        when x"13D7" => data_out<= x"20";
        when x"13D8" => data_out<= x"93";
        when x"13D9" => data_out<= x"B0";
        when x"13DA" => data_out<= x"A9";
        when x"13DB" => data_out<= x"0A";
        when x"13DC" => data_out<= x"20";
        when x"13DD" => data_out<= x"20";
        when x"13DE" => data_out<= x"B1";
        when x"13DF" => data_out<= x"A0";
        when x"13E0" => data_out<= x"07";
        when x"13E1" => data_out<= x"20";
        when x"13E2" => data_out<= x"C5";
        when x"13E3" => data_out<= x"B0";
        when x"13E4" => data_out<= x"A0";
        when x"13E5" => data_out<= x"07";
        when x"13E6" => data_out<= x"B1";
        when x"13E7" => data_out<= x"0C";
        when x"13E8" => data_out<= x"C8";
        when x"13E9" => data_out<= x"11";
        when x"13EA" => data_out<= x"0C";
        when x"13EB" => data_out<= x"D0";
        when x"13EC" => data_out<= x"B5";
        when x"13ED" => data_out<= x"4C";
        when x"13EE" => data_out<= x"0F";
        when x"13EF" => data_out<= x"94";
        when x"13F0" => data_out<= x"B1";
        when x"13F1" => data_out<= x"0C";
        when x"13F2" => data_out<= x"38";
        when x"13F3" => data_out<= x"E9";
        when x"13F4" => data_out<= x"01";
        when x"13F5" => data_out<= x"91";
        when x"13F6" => data_out<= x"0C";
        when x"13F7" => data_out<= x"18";
        when x"13F8" => data_out<= x"69";
        when x"13F9" => data_out<= x"01";
        when x"13FA" => data_out<= x"90";
        when x"13FB" => data_out<= x"03";
        when x"13FC" => data_out<= x"A2";
        when x"13FD" => data_out<= x"01";
        when x"13FE" => data_out<= x"18";
        when x"13FF" => data_out<= x"65";
        when x"1400" => data_out<= x"0C";
        when x"1401" => data_out<= x"85";
        when x"1402" => data_out<= x"14";
        when x"1403" => data_out<= x"8A";
        when x"1404" => data_out<= x"65";
        when x"1405" => data_out<= x"0D";
        when x"1406" => data_out<= x"85";
        when x"1407" => data_out<= x"15";
        when x"1408" => data_out<= x"A0";
        when x"1409" => data_out<= x"00";
        when x"140A" => data_out<= x"B1";
        when x"140B" => data_out<= x"14";
        when x"140C" => data_out<= x"20";
        when x"140D" => data_out<= x"F0";
        when x"140E" => data_out<= x"80";
        when x"140F" => data_out<= x"A0";
        when x"1410" => data_out<= x"00";
        when x"1411" => data_out<= x"A2";
        when x"1412" => data_out<= x"00";
        when x"1413" => data_out<= x"B1";
        when x"1414" => data_out<= x"0C";
        when x"1415" => data_out<= x"D0";
        when x"1416" => data_out<= x"D9";
        when x"1417" => data_out<= x"A0";
        when x"1418" => data_out<= x"09";
        when x"1419" => data_out<= x"4C";
        when x"141A" => data_out<= x"14";
        when x"141B" => data_out<= x"AE";
        when x"141C" => data_out<= x"20";
        when x"141D" => data_out<= x"45";
        when x"141E" => data_out<= x"8C";
        when x"141F" => data_out<= x"A9";
        when x"1420" => data_out<= x"9E";
        when x"1421" => data_out<= x"A2";
        when x"1422" => data_out<= x"B8";
        when x"1423" => data_out<= x"20";
        when x"1424" => data_out<= x"22";
        when x"1425" => data_out<= x"81";
        when x"1426" => data_out<= x"20";
        when x"1427" => data_out<= x"45";
        when x"1428" => data_out<= x"8C";
        when x"1429" => data_out<= x"20";
        when x"142A" => data_out<= x"45";
        when x"142B" => data_out<= x"8C";
        when x"142C" => data_out<= x"A9";
        when x"142D" => data_out<= x"FA";
        when x"142E" => data_out<= x"A2";
        when x"142F" => data_out<= x"B6";
        when x"1430" => data_out<= x"20";
        when x"1431" => data_out<= x"22";
        when x"1432" => data_out<= x"81";
        when x"1433" => data_out<= x"A2";
        when x"1434" => data_out<= x"00";
        when x"1435" => data_out<= x"A9";
        when x"1436" => data_out<= x"FE";
        when x"1437" => data_out<= x"20";
        when x"1438" => data_out<= x"86";
        when x"1439" => data_out<= x"93";
        when x"143A" => data_out<= x"A9";
        when x"143B" => data_out<= x"1C";
        when x"143C" => data_out<= x"A2";
        when x"143D" => data_out<= x"BC";
        when x"143E" => data_out<= x"20";
        when x"143F" => data_out<= x"22";
        when x"1440" => data_out<= x"81";
        when x"1441" => data_out<= x"20";
        when x"1442" => data_out<= x"45";
        when x"1443" => data_out<= x"8C";
        when x"1444" => data_out<= x"A9";
        when x"1445" => data_out<= x"E0";
        when x"1446" => data_out<= x"A2";
        when x"1447" => data_out<= x"B6";
        when x"1448" => data_out<= x"20";
        when x"1449" => data_out<= x"22";
        when x"144A" => data_out<= x"81";
        when x"144B" => data_out<= x"A2";
        when x"144C" => data_out<= x"3D";
        when x"144D" => data_out<= x"A9";
        when x"144E" => data_out<= x"00";
        when x"144F" => data_out<= x"20";
        when x"1450" => data_out<= x"86";
        when x"1451" => data_out<= x"93";
        when x"1452" => data_out<= x"A9";
        when x"1453" => data_out<= x"1C";
        when x"1454" => data_out<= x"A2";
        when x"1455" => data_out<= x"BC";
        when x"1456" => data_out<= x"20";
        when x"1457" => data_out<= x"22";
        when x"1458" => data_out<= x"81";
        when x"1459" => data_out<= x"20";
        when x"145A" => data_out<= x"45";
        when x"145B" => data_out<= x"8C";
        when x"145C" => data_out<= x"A9";
        when x"145D" => data_out<= x"2E";
        when x"145E" => data_out<= x"A2";
        when x"145F" => data_out<= x"B7";
        when x"1460" => data_out<= x"20";
        when x"1461" => data_out<= x"22";
        when x"1462" => data_out<= x"81";
        when x"1463" => data_out<= x"A2";
        when x"1464" => data_out<= x"02";
        when x"1465" => data_out<= x"A9";
        when x"1466" => data_out<= x"00";
        when x"1467" => data_out<= x"20";
        when x"1468" => data_out<= x"86";
        when x"1469" => data_out<= x"93";
        when x"146A" => data_out<= x"A9";
        when x"146B" => data_out<= x"1C";
        when x"146C" => data_out<= x"A2";
        when x"146D" => data_out<= x"BC";
        when x"146E" => data_out<= x"20";
        when x"146F" => data_out<= x"22";
        when x"1470" => data_out<= x"81";
        when x"1471" => data_out<= x"20";
        when x"1472" => data_out<= x"45";
        when x"1473" => data_out<= x"8C";
        when x"1474" => data_out<= x"A9";
        when x"1475" => data_out<= x"F5";
        when x"1476" => data_out<= x"A2";
        when x"1477" => data_out<= x"B3";
        when x"1478" => data_out<= x"20";
        when x"1479" => data_out<= x"22";
        when x"147A" => data_out<= x"81";
        when x"147B" => data_out<= x"20";
        when x"147C" => data_out<= x"45";
        when x"147D" => data_out<= x"8C";
        when x"147E" => data_out<= x"A9";
        when x"147F" => data_out<= x"C6";
        when x"1480" => data_out<= x"A2";
        when x"1481" => data_out<= x"B7";
        when x"1482" => data_out<= x"20";
        when x"1483" => data_out<= x"22";
        when x"1484" => data_out<= x"81";
        when x"1485" => data_out<= x"20";
        when x"1486" => data_out<= x"45";
        when x"1487" => data_out<= x"8C";
        when x"1488" => data_out<= x"20";
        when x"1489" => data_out<= x"45";
        when x"148A" => data_out<= x"8C";
        when x"148B" => data_out<= x"A9";
        when x"148C" => data_out<= x"95";
        when x"148D" => data_out<= x"A2";
        when x"148E" => data_out<= x"B7";
        when x"148F" => data_out<= x"20";
        when x"1490" => data_out<= x"22";
        when x"1491" => data_out<= x"81";
        when x"1492" => data_out<= x"20";
        when x"1493" => data_out<= x"45";
        when x"1494" => data_out<= x"8C";
        when x"1495" => data_out<= x"A9";
        when x"1496" => data_out<= x"E8";
        when x"1497" => data_out<= x"A2";
        when x"1498" => data_out<= x"B9";
        when x"1499" => data_out<= x"20";
        when x"149A" => data_out<= x"22";
        when x"149B" => data_out<= x"81";
        when x"149C" => data_out<= x"20";
        when x"149D" => data_out<= x"45";
        when x"149E" => data_out<= x"8C";
        when x"149F" => data_out<= x"A9";
        when x"14A0" => data_out<= x"27";
        when x"14A1" => data_out<= x"A2";
        when x"14A2" => data_out<= x"BB";
        when x"14A3" => data_out<= x"20";
        when x"14A4" => data_out<= x"22";
        when x"14A5" => data_out<= x"81";
        when x"14A6" => data_out<= x"A2";
        when x"14A7" => data_out<= x"36";
        when x"14A8" => data_out<= x"A9";
        when x"14A9" => data_out<= x"00";
        when x"14AA" => data_out<= x"20";
        when x"14AB" => data_out<= x"86";
        when x"14AC" => data_out<= x"93";
        when x"14AD" => data_out<= x"A9";
        when x"14AE" => data_out<= x"1C";
        when x"14AF" => data_out<= x"A2";
        when x"14B0" => data_out<= x"BC";
        when x"14B1" => data_out<= x"20";
        when x"14B2" => data_out<= x"22";
        when x"14B3" => data_out<= x"81";
        when x"14B4" => data_out<= x"4C";
        when x"14B5" => data_out<= x"45";
        when x"14B6" => data_out<= x"8C";
        when x"14B7" => data_out<= x"20";
        when x"14B8" => data_out<= x"6A";
        when x"14B9" => data_out<= x"AE";
        when x"14BA" => data_out<= x"A9";
        when x"14BB" => data_out<= x"7C";
        when x"14BC" => data_out<= x"A2";
        when x"14BD" => data_out<= x"B7";
        when x"14BE" => data_out<= x"20";
        when x"14BF" => data_out<= x"22";
        when x"14C0" => data_out<= x"81";
        when x"14C1" => data_out<= x"20";
        when x"14C2" => data_out<= x"45";
        when x"14C3" => data_out<= x"8C";
        when x"14C4" => data_out<= x"20";
        when x"14C5" => data_out<= x"BF";
        when x"14C6" => data_out<= x"9F";
        when x"14C7" => data_out<= x"A0";
        when x"14C8" => data_out<= x"00";
        when x"14C9" => data_out<= x"91";
        when x"14CA" => data_out<= x"0C";
        when x"14CB" => data_out<= x"B1";
        when x"14CC" => data_out<= x"0C";
        when x"14CD" => data_out<= x"F0";
        when x"14CE" => data_out<= x"1C";
        when x"14CF" => data_out<= x"A9";
        when x"14D0" => data_out<= x"A4";
        when x"14D1" => data_out<= x"A2";
        when x"14D2" => data_out<= x"BB";
        when x"14D3" => data_out<= x"20";
        when x"14D4" => data_out<= x"22";
        when x"14D5" => data_out<= x"81";
        when x"14D6" => data_out<= x"A0";
        when x"14D7" => data_out<= x"00";
        when x"14D8" => data_out<= x"B1";
        when x"14D9" => data_out<= x"0C";
        when x"14DA" => data_out<= x"20";
        when x"14DB" => data_out<= x"FD";
        when x"14DC" => data_out<= x"8B";
        when x"14DD" => data_out<= x"20";
        when x"14DE" => data_out<= x"45";
        when x"14DF" => data_out<= x"8C";
        when x"14E0" => data_out<= x"A9";
        when x"14E1" => data_out<= x"00";
        when x"14E2" => data_out<= x"8D";
        when x"14E3" => data_out<= x"02";
        when x"14E4" => data_out<= x"02";
        when x"14E5" => data_out<= x"8D";
        when x"14E6" => data_out<= x"03";
        when x"14E7" => data_out<= x"02";
        when x"14E8" => data_out<= x"4C";
        when x"14E9" => data_out<= x"05";
        when x"14EA" => data_out<= x"AF";
        when x"14EB" => data_out<= x"A9";
        when x"14EC" => data_out<= x"01";
        when x"14ED" => data_out<= x"8D";
        when x"14EE" => data_out<= x"02";
        when x"14EF" => data_out<= x"02";
        when x"14F0" => data_out<= x"A9";
        when x"14F1" => data_out<= x"B7";
        when x"14F2" => data_out<= x"A2";
        when x"14F3" => data_out<= x"BA";
        when x"14F4" => data_out<= x"20";
        when x"14F5" => data_out<= x"22";
        when x"14F6" => data_out<= x"81";
        when x"14F7" => data_out<= x"20";
        when x"14F8" => data_out<= x"71";
        when x"14F9" => data_out<= x"A2";
        when x"14FA" => data_out<= x"C9";
        when x"14FB" => data_out<= x"02";
        when x"14FC" => data_out<= x"D0";
        when x"14FD" => data_out<= x"05";
        when x"14FE" => data_out<= x"A9";
        when x"14FF" => data_out<= x"48";
        when x"1500" => data_out<= x"4C";
        when x"1501" => data_out<= x"05";
        when x"1502" => data_out<= x"95";
        when x"1503" => data_out<= x"A9";
        when x"1504" => data_out<= x"53";
        when x"1505" => data_out<= x"20";
        when x"1506" => data_out<= x"F0";
        when x"1507" => data_out<= x"80";
        when x"1508" => data_out<= x"A9";
        when x"1509" => data_out<= x"44";
        when x"150A" => data_out<= x"20";
        when x"150B" => data_out<= x"F0";
        when x"150C" => data_out<= x"80";
        when x"150D" => data_out<= x"20";
        when x"150E" => data_out<= x"45";
        when x"150F" => data_out<= x"8C";
        when x"1510" => data_out<= x"A9";
        when x"1511" => data_out<= x"FC";
        when x"1512" => data_out<= x"A2";
        when x"1513" => data_out<= x"B9";
        when x"1514" => data_out<= x"20";
        when x"1515" => data_out<= x"22";
        when x"1516" => data_out<= x"81";
        when x"1517" => data_out<= x"20";
        when x"1518" => data_out<= x"45";
        when x"1519" => data_out<= x"8C";
        when x"151A" => data_out<= x"20";
        when x"151B" => data_out<= x"68";
        when x"151C" => data_out<= x"A3";
        when x"151D" => data_out<= x"A0";
        when x"151E" => data_out<= x"00";
        when x"151F" => data_out<= x"91";
        when x"1520" => data_out<= x"0C";
        when x"1521" => data_out<= x"C9";
        when x"1522" => data_out<= x"02";
        when x"1523" => data_out<= x"D0";
        when x"1524" => data_out<= x"3B";
        when x"1525" => data_out<= x"A9";
        when x"1526" => data_out<= x"7F";
        when x"1527" => data_out<= x"A2";
        when x"1528" => data_out<= x"B5";
        when x"1529" => data_out<= x"20";
        when x"152A" => data_out<= x"22";
        when x"152B" => data_out<= x"81";
        when x"152C" => data_out<= x"20";
        when x"152D" => data_out<= x"FD";
        when x"152E" => data_out<= x"80";
        when x"152F" => data_out<= x"C9";
        when x"1530" => data_out<= x"53";
        when x"1531" => data_out<= x"F0";
        when x"1532" => data_out<= x"07";
        when x"1533" => data_out<= x"20";
        when x"1534" => data_out<= x"FD";
        when x"1535" => data_out<= x"80";
        when x"1536" => data_out<= x"C9";
        when x"1537" => data_out<= x"73";
        when x"1538" => data_out<= x"D0";
        when x"1539" => data_out<= x"47";
        when x"153A" => data_out<= x"20";
        when x"153B" => data_out<= x"45";
        when x"153C" => data_out<= x"8C";
        when x"153D" => data_out<= x"A9";
        when x"153E" => data_out<= x"A6";
        when x"153F" => data_out<= x"A2";
        when x"1540" => data_out<= x"BA";
        when x"1541" => data_out<= x"20";
        when x"1542" => data_out<= x"22";
        when x"1543" => data_out<= x"81";
        when x"1544" => data_out<= x"20";
        when x"1545" => data_out<= x"9D";
        when x"1546" => data_out<= x"A3";
        when x"1547" => data_out<= x"A0";
        when x"1548" => data_out<= x"00";
        when x"1549" => data_out<= x"91";
        when x"154A" => data_out<= x"0C";
        when x"154B" => data_out<= x"B1";
        when x"154C" => data_out<= x"0C";
        when x"154D" => data_out<= x"D0";
        when x"154E" => data_out<= x"11";
        when x"154F" => data_out<= x"A9";
        when x"1550" => data_out<= x"F4";
        when x"1551" => data_out<= x"A2";
        when x"1552" => data_out<= x"BA";
        when x"1553" => data_out<= x"20";
        when x"1554" => data_out<= x"22";
        when x"1555" => data_out<= x"81";
        when x"1556" => data_out<= x"20";
        when x"1557" => data_out<= x"45";
        when x"1558" => data_out<= x"8C";
        when x"1559" => data_out<= x"20";
        when x"155A" => data_out<= x"68";
        when x"155B" => data_out<= x"A3";
        when x"155C" => data_out<= x"A0";
        when x"155D" => data_out<= x"00";
        when x"155E" => data_out<= x"91";
        when x"155F" => data_out<= x"0C";
        when x"1560" => data_out<= x"B1";
        when x"1561" => data_out<= x"0C";
        when x"1562" => data_out<= x"D0";
        when x"1563" => data_out<= x"0F";
        when x"1564" => data_out<= x"A9";
        when x"1565" => data_out<= x"01";
        when x"1566" => data_out<= x"8D";
        when x"1567" => data_out<= x"03";
        when x"1568" => data_out<= x"02";
        when x"1569" => data_out<= x"A9";
        when x"156A" => data_out<= x"E7";
        when x"156B" => data_out<= x"A2";
        when x"156C" => data_out<= x"BA";
        when x"156D" => data_out<= x"20";
        when x"156E" => data_out<= x"22";
        when x"156F" => data_out<= x"81";
        when x"1570" => data_out<= x"4C";
        when x"1571" => data_out<= x"81";
        when x"1572" => data_out<= x"95";
        when x"1573" => data_out<= x"A9";
        when x"1574" => data_out<= x"B1";
        when x"1575" => data_out<= x"A2";
        when x"1576" => data_out<= x"BB";
        when x"1577" => data_out<= x"20";
        when x"1578" => data_out<= x"22";
        when x"1579" => data_out<= x"81";
        when x"157A" => data_out<= x"A0";
        when x"157B" => data_out<= x"00";
        when x"157C" => data_out<= x"B1";
        when x"157D" => data_out<= x"0C";
        when x"157E" => data_out<= x"20";
        when x"157F" => data_out<= x"FD";
        when x"1580" => data_out<= x"8B";
        when x"1581" => data_out<= x"20";
        when x"1582" => data_out<= x"45";
        when x"1583" => data_out<= x"8C";
        when x"1584" => data_out<= x"4C";
        when x"1585" => data_out<= x"05";
        when x"1586" => data_out<= x"AF";
        when x"1587" => data_out<= x"A0";
        when x"1588" => data_out<= x"10";
        when x"1589" => data_out<= x"20";
        when x"158A" => data_out<= x"13";
        when x"158B" => data_out<= x"B1";
        when x"158C" => data_out<= x"A9";
        when x"158D" => data_out<= x"00";
        when x"158E" => data_out<= x"20";
        when x"158F" => data_out<= x"65";
        when x"1590" => data_out<= x"B0";
        when x"1591" => data_out<= x"AD";
        when x"1592" => data_out<= x"03";
        when x"1593" => data_out<= x"02";
        when x"1594" => data_out<= x"D0";
        when x"1595" => data_out<= x"07";
        when x"1596" => data_out<= x"A9";
        when x"1597" => data_out<= x"B1";
        when x"1598" => data_out<= x"A2";
        when x"1599" => data_out<= x"B4";
        when x"159A" => data_out<= x"4C";
        when x"159B" => data_out<= x"20";
        when x"159C" => data_out<= x"96";
        when x"159D" => data_out<= x"A9";
        when x"159E" => data_out<= x"00";
        when x"159F" => data_out<= x"A2";
        when x"15A0" => data_out<= x"BC";
        when x"15A1" => data_out<= x"20";
        when x"15A2" => data_out<= x"22";
        when x"15A3" => data_out<= x"81";
        when x"15A4" => data_out<= x"20";
        when x"15A5" => data_out<= x"45";
        when x"15A6" => data_out<= x"8C";
        when x"15A7" => data_out<= x"A9";
        when x"15A8" => data_out<= x"00";
        when x"15A9" => data_out<= x"A0";
        when x"15AA" => data_out<= x"01";
        when x"15AB" => data_out<= x"91";
        when x"15AC" => data_out<= x"0C";
        when x"15AD" => data_out<= x"C9";
        when x"15AE" => data_out<= x"10";
        when x"15AF" => data_out<= x"B0";
        when x"15B0" => data_out<= x"4C";
        when x"15B1" => data_out<= x"B1";
        when x"15B2" => data_out<= x"0C";
        when x"15B3" => data_out<= x"20";
        when x"15B4" => data_out<= x"65";
        when x"15B5" => data_out<= x"B0";
        when x"15B6" => data_out<= x"A9";
        when x"15B7" => data_out<= x"03";
        when x"15B8" => data_out<= x"20";
        when x"15B9" => data_out<= x"69";
        when x"15BA" => data_out<= x"AF";
        when x"15BB" => data_out<= x"20";
        when x"15BC" => data_out<= x"51";
        when x"15BD" => data_out<= x"AA";
        when x"15BE" => data_out<= x"C9";
        when x"15BF" => data_out<= x"00";
        when x"15C0" => data_out<= x"D0";
        when x"15C1" => data_out<= x"31";
        when x"15C2" => data_out<= x"A9";
        when x"15C3" => data_out<= x"02";
        when x"15C4" => data_out<= x"A2";
        when x"15C5" => data_out<= x"BD";
        when x"15C6" => data_out<= x"20";
        when x"15C7" => data_out<= x"22";
        when x"15C8" => data_out<= x"81";
        when x"15C9" => data_out<= x"A9";
        when x"15CA" => data_out<= x"02";
        when x"15CB" => data_out<= x"20";
        when x"15CC" => data_out<= x"69";
        when x"15CD" => data_out<= x"AF";
        when x"15CE" => data_out<= x"20";
        when x"15CF" => data_out<= x"22";
        when x"15D0" => data_out<= x"81";
        when x"15D1" => data_out<= x"A9";
        when x"15D2" => data_out<= x"02";
        when x"15D3" => data_out<= x"A2";
        when x"15D4" => data_out<= x"BD";
        when x"15D5" => data_out<= x"20";
        when x"15D6" => data_out<= x"22";
        when x"15D7" => data_out<= x"81";
        when x"15D8" => data_out<= x"A0";
        when x"15D9" => data_out<= x"0F";
        when x"15DA" => data_out<= x"20";
        when x"15DB" => data_out<= x"4F";
        when x"15DC" => data_out<= x"AF";
        when x"15DD" => data_out<= x"20";
        when x"15DE" => data_out<= x"86";
        when x"15DF" => data_out<= x"93";
        when x"15E0" => data_out<= x"A9";
        when x"15E1" => data_out<= x"34";
        when x"15E2" => data_out<= x"A2";
        when x"15E3" => data_out<= x"BC";
        when x"15E4" => data_out<= x"20";
        when x"15E5" => data_out<= x"22";
        when x"15E6" => data_out<= x"81";
        when x"15E7" => data_out<= x"20";
        when x"15E8" => data_out<= x"45";
        when x"15E9" => data_out<= x"8C";
        when x"15EA" => data_out<= x"A0";
        when x"15EB" => data_out<= x"00";
        when x"15EC" => data_out<= x"B1";
        when x"15ED" => data_out<= x"0C";
        when x"15EE" => data_out<= x"18";
        when x"15EF" => data_out<= x"69";
        when x"15F0" => data_out<= x"01";
        when x"15F1" => data_out<= x"91";
        when x"15F2" => data_out<= x"0C";
        when x"15F3" => data_out<= x"A0";
        when x"15F4" => data_out<= x"01";
        when x"15F5" => data_out<= x"B1";
        when x"15F6" => data_out<= x"0C";
        when x"15F7" => data_out<= x"18";
        when x"15F8" => data_out<= x"69";
        when x"15F9" => data_out<= x"01";
        when x"15FA" => data_out<= x"4C";
        when x"15FB" => data_out<= x"AB";
        when x"15FC" => data_out<= x"95";
        when x"15FD" => data_out<= x"88";
        when x"15FE" => data_out<= x"B1";
        when x"15FF" => data_out<= x"0C";
        when x"1600" => data_out<= x"D0";
        when x"1601" => data_out<= x"0A";
        when x"1602" => data_out<= x"A9";
        when x"1603" => data_out<= x"F6";
        when x"1604" => data_out<= x"A2";
        when x"1605" => data_out<= x"BB";
        when x"1606" => data_out<= x"20";
        when x"1607" => data_out<= x"22";
        when x"1608" => data_out<= x"81";
        when x"1609" => data_out<= x"20";
        when x"160A" => data_out<= x"45";
        when x"160B" => data_out<= x"8C";
        when x"160C" => data_out<= x"A9";
        when x"160D" => data_out<= x"24";
        when x"160E" => data_out<= x"A2";
        when x"160F" => data_out<= x"BC";
        when x"1610" => data_out<= x"20";
        when x"1611" => data_out<= x"22";
        when x"1612" => data_out<= x"81";
        when x"1613" => data_out<= x"A0";
        when x"1614" => data_out<= x"00";
        when x"1615" => data_out<= x"B1";
        when x"1616" => data_out<= x"0C";
        when x"1617" => data_out<= x"A2";
        when x"1618" => data_out<= x"00";
        when x"1619" => data_out<= x"20";
        when x"161A" => data_out<= x"86";
        when x"161B" => data_out<= x"93";
        when x"161C" => data_out<= x"A9";
        when x"161D" => data_out<= x"70";
        when x"161E" => data_out<= x"A2";
        when x"161F" => data_out<= x"BB";
        when x"1620" => data_out<= x"20";
        when x"1621" => data_out<= x"22";
        when x"1622" => data_out<= x"81";
        when x"1623" => data_out<= x"20";
        when x"1624" => data_out<= x"45";
        when x"1625" => data_out<= x"8C";
        when x"1626" => data_out<= x"A0";
        when x"1627" => data_out<= x"11";
        when x"1628" => data_out<= x"4C";
        when x"1629" => data_out<= x"14";
        when x"162A" => data_out<= x"AE";
        when x"162B" => data_out<= x"20";
        when x"162C" => data_out<= x"7B";
        when x"162D" => data_out<= x"B0";
        when x"162E" => data_out<= x"20";
        when x"162F" => data_out<= x"6A";
        when x"1630" => data_out<= x"AE";
        when x"1631" => data_out<= x"20";
        when x"1632" => data_out<= x"77";
        when x"1633" => data_out<= x"B0";
        when x"1634" => data_out<= x"A0";
        when x"1635" => data_out<= x"44";
        when x"1636" => data_out<= x"20";
        when x"1637" => data_out<= x"13";
        when x"1638" => data_out<= x"B1";
        when x"1639" => data_out<= x"AD";
        when x"163A" => data_out<= x"03";
        when x"163B" => data_out<= x"02";
        when x"163C" => data_out<= x"D0";
        when x"163D" => data_out<= x"07";
        when x"163E" => data_out<= x"A9";
        when x"163F" => data_out<= x"46";
        when x"1640" => data_out<= x"A2";
        when x"1641" => data_out<= x"BB";
        when x"1642" => data_out<= x"4C";
        when x"1643" => data_out<= x"A4";
        when x"1644" => data_out<= x"97";
        when x"1645" => data_out<= x"A0";
        when x"1646" => data_out<= x"47";
        when x"1647" => data_out<= x"B1";
        when x"1648" => data_out<= x"0C";
        when x"1649" => data_out<= x"C8";
        when x"164A" => data_out<= x"11";
        when x"164B" => data_out<= x"0C";
        when x"164C" => data_out<= x"F0";
        when x"164D" => data_out<= x"0A";
        when x"164E" => data_out<= x"20";
        when x"164F" => data_out<= x"4F";
        when x"1650" => data_out<= x"AF";
        when x"1651" => data_out<= x"C9";
        when x"1652" => data_out<= x"01";
        when x"1653" => data_out<= x"8A";
        when x"1654" => data_out<= x"E9";
        when x"1655" => data_out<= x"80";
        when x"1656" => data_out<= x"90";
        when x"1657" => data_out<= x"07";
        when x"1658" => data_out<= x"A9";
        when x"1659" => data_out<= x"12";
        when x"165A" => data_out<= x"A2";
        when x"165B" => data_out<= x"B9";
        when x"165C" => data_out<= x"4C";
        when x"165D" => data_out<= x"A4";
        when x"165E" => data_out<= x"97";
        when x"165F" => data_out<= x"A0";
        when x"1660" => data_out<= x"4C";
        when x"1661" => data_out<= x"20";
        when x"1662" => data_out<= x"4F";
        when x"1663" => data_out<= x"AF";
        when x"1664" => data_out<= x"20";
        when x"1665" => data_out<= x"DF";
        when x"1666" => data_out<= x"A9";
        when x"1667" => data_out<= x"A0";
        when x"1668" => data_out<= x"4E";
        when x"1669" => data_out<= x"20";
        when x"166A" => data_out<= x"93";
        when x"166B" => data_out<= x"B0";
        when x"166C" => data_out<= x"A0";
        when x"166D" => data_out<= x"4A";
        when x"166E" => data_out<= x"20";
        when x"166F" => data_out<= x"4F";
        when x"1670" => data_out<= x"AF";
        when x"1671" => data_out<= x"20";
        when x"1672" => data_out<= x"BC";
        when x"1673" => data_out<= x"A4";
        when x"1674" => data_out<= x"A0";
        when x"1675" => data_out<= x"46";
        when x"1676" => data_out<= x"91";
        when x"1677" => data_out<= x"0C";
        when x"1678" => data_out<= x"B1";
        when x"1679" => data_out<= x"0C";
        when x"167A" => data_out<= x"F0";
        when x"167B" => data_out<= x"11";
        when x"167C" => data_out<= x"A9";
        when x"167D" => data_out<= x"62";
        when x"167E" => data_out<= x"A2";
        when x"167F" => data_out<= x"BB";
        when x"1680" => data_out<= x"20";
        when x"1681" => data_out<= x"22";
        when x"1682" => data_out<= x"81";
        when x"1683" => data_out<= x"A0";
        when x"1684" => data_out<= x"46";
        when x"1685" => data_out<= x"B1";
        when x"1686" => data_out<= x"0C";
        when x"1687" => data_out<= x"20";
        when x"1688" => data_out<= x"FD";
        when x"1689" => data_out<= x"8B";
        when x"168A" => data_out<= x"4C";
        when x"168B" => data_out<= x"A7";
        when x"168C" => data_out<= x"97";
        when x"168D" => data_out<= x"A9";
        when x"168E" => data_out<= x"BE";
        when x"168F" => data_out<= x"A2";
        when x"1690" => data_out<= x"BB";
        when x"1691" => data_out<= x"20";
        when x"1692" => data_out<= x"22";
        when x"1693" => data_out<= x"81";
        when x"1694" => data_out<= x"A0";
        when x"1695" => data_out<= x"4A";
        when x"1696" => data_out<= x"20";
        when x"1697" => data_out<= x"4F";
        when x"1698" => data_out<= x"AF";
        when x"1699" => data_out<= x"20";
        when x"169A" => data_out<= x"31";
        when x"169B" => data_out<= x"8C";
        when x"169C" => data_out<= x"A9";
        when x"169D" => data_out<= x"7D";
        when x"169E" => data_out<= x"A2";
        when x"169F" => data_out<= x"BD";
        when x"16A0" => data_out<= x"20";
        when x"16A1" => data_out<= x"22";
        when x"16A2" => data_out<= x"81";
        when x"16A3" => data_out<= x"A0";
        when x"16A4" => data_out<= x"48";
        when x"16A5" => data_out<= x"20";
        when x"16A6" => data_out<= x"4F";
        when x"16A7" => data_out<= x"AF";
        when x"16A8" => data_out<= x"18";
        when x"16A9" => data_out<= x"A0";
        when x"16AA" => data_out<= x"49";
        when x"16AB" => data_out<= x"71";
        when x"16AC" => data_out<= x"0C";
        when x"16AD" => data_out<= x"48";
        when x"16AE" => data_out<= x"8A";
        when x"16AF" => data_out<= x"C8";
        when x"16B0" => data_out<= x"71";
        when x"16B1" => data_out<= x"0C";
        when x"16B2" => data_out<= x"AA";
        when x"16B3" => data_out<= x"68";
        when x"16B4" => data_out<= x"20";
        when x"16B5" => data_out<= x"5A";
        when x"16B6" => data_out<= x"AE";
        when x"16B7" => data_out<= x"20";
        when x"16B8" => data_out<= x"31";
        when x"16B9" => data_out<= x"8C";
        when x"16BA" => data_out<= x"A9";
        when x"16BB" => data_out<= x"8B";
        when x"16BC" => data_out<= x"A2";
        when x"16BD" => data_out<= x"BC";
        when x"16BE" => data_out<= x"20";
        when x"16BF" => data_out<= x"22";
        when x"16C0" => data_out<= x"81";
        when x"16C1" => data_out<= x"A0";
        when x"16C2" => data_out<= x"4C";
        when x"16C3" => data_out<= x"20";
        when x"16C4" => data_out<= x"4F";
        when x"16C5" => data_out<= x"AF";
        when x"16C6" => data_out<= x"20";
        when x"16C7" => data_out<= x"22";
        when x"16C8" => data_out<= x"81";
        when x"16C9" => data_out<= x"20";
        when x"16CA" => data_out<= x"45";
        when x"16CB" => data_out<= x"8C";
        when x"16CC" => data_out<= x"4C";
        when x"16CD" => data_out<= x"79";
        when x"16CE" => data_out<= x"97";
        when x"16CF" => data_out<= x"20";
        when x"16D0" => data_out<= x"4F";
        when x"16D1" => data_out<= x"AF";
        when x"16D2" => data_out<= x"38";
        when x"16D3" => data_out<= x"A0";
        when x"16D4" => data_out<= x"44";
        when x"16D5" => data_out<= x"F1";
        when x"16D6" => data_out<= x"0C";
        when x"16D7" => data_out<= x"48";
        when x"16D8" => data_out<= x"8A";
        when x"16D9" => data_out<= x"C8";
        when x"16DA" => data_out<= x"F1";
        when x"16DB" => data_out<= x"0C";
        when x"16DC" => data_out<= x"AA";
        when x"16DD" => data_out<= x"68";
        when x"16DE" => data_out<= x"A0";
        when x"16DF" => data_out<= x"42";
        when x"16E0" => data_out<= x"20";
        when x"16E1" => data_out<= x"C5";
        when x"16E2" => data_out<= x"B0";
        when x"16E3" => data_out<= x"C9";
        when x"16E4" => data_out<= x"41";
        when x"16E5" => data_out<= x"8A";
        when x"16E6" => data_out<= x"E9";
        when x"16E7" => data_out<= x"00";
        when x"16E8" => data_out<= x"A9";
        when x"16E9" => data_out<= x"00";
        when x"16EA" => data_out<= x"AA";
        when x"16EB" => data_out<= x"90";
        when x"16EC" => data_out<= x"08";
        when x"16ED" => data_out<= x"A9";
        when x"16EE" => data_out<= x"40";
        when x"16EF" => data_out<= x"A0";
        when x"16F0" => data_out<= x"42";
        when x"16F1" => data_out<= x"20";
        when x"16F2" => data_out<= x"C5";
        when x"16F3" => data_out<= x"B0";
        when x"16F4" => data_out<= x"8A";
        when x"16F5" => data_out<= x"20";
        when x"16F6" => data_out<= x"C3";
        when x"16F7" => data_out<= x"B0";
        when x"16F8" => data_out<= x"A0";
        when x"16F9" => data_out<= x"42";
        when x"16FA" => data_out<= x"D1";
        when x"16FB" => data_out<= x"0C";
        when x"16FC" => data_out<= x"8A";
        when x"16FD" => data_out<= x"C8";
        when x"16FE" => data_out<= x"F1";
        when x"16FF" => data_out<= x"0C";
        when x"1700" => data_out<= x"B0";
        when x"1701" => data_out<= x"45";
        when x"1702" => data_out<= x"A9";
        when x"1703" => data_out<= x"02";
        when x"1704" => data_out<= x"20";
        when x"1705" => data_out<= x"69";
        when x"1706" => data_out<= x"AF";
        when x"1707" => data_out<= x"A0";
        when x"1708" => data_out<= x"00";
        when x"1709" => data_out<= x"18";
        when x"170A" => data_out<= x"71";
        when x"170B" => data_out<= x"0C";
        when x"170C" => data_out<= x"48";
        when x"170D" => data_out<= x"8A";
        when x"170E" => data_out<= x"C8";
        when x"170F" => data_out<= x"71";
        when x"1710" => data_out<= x"0C";
        when x"1711" => data_out<= x"AA";
        when x"1712" => data_out<= x"68";
        when x"1713" => data_out<= x"20";
        when x"1714" => data_out<= x"7B";
        when x"1715" => data_out<= x"B0";
        when x"1716" => data_out<= x"A0";
        when x"1717" => data_out<= x"47";
        when x"1718" => data_out<= x"20";
        when x"1719" => data_out<= x"4F";
        when x"171A" => data_out<= x"AF";
        when x"171B" => data_out<= x"18";
        when x"171C" => data_out<= x"A0";
        when x"171D" => data_out<= x"4B";
        when x"171E" => data_out<= x"71";
        when x"171F" => data_out<= x"0C";
        when x"1720" => data_out<= x"85";
        when x"1721" => data_out<= x"14";
        when x"1722" => data_out<= x"8A";
        when x"1723" => data_out<= x"C8";
        when x"1724" => data_out<= x"71";
        when x"1725" => data_out<= x"0C";
        when x"1726" => data_out<= x"85";
        when x"1727" => data_out<= x"15";
        when x"1728" => data_out<= x"A0";
        when x"1729" => data_out<= x"03";
        when x"172A" => data_out<= x"20";
        when x"172B" => data_out<= x"4F";
        when x"172C" => data_out<= x"AF";
        when x"172D" => data_out<= x"18";
        when x"172E" => data_out<= x"65";
        when x"172F" => data_out<= x"14";
        when x"1730" => data_out<= x"48";
        when x"1731" => data_out<= x"8A";
        when x"1732" => data_out<= x"65";
        when x"1733" => data_out<= x"15";
        when x"1734" => data_out<= x"AA";
        when x"1735" => data_out<= x"68";
        when x"1736" => data_out<= x"20";
        when x"1737" => data_out<= x"49";
        when x"1738" => data_out<= x"89";
        when x"1739" => data_out<= x"A0";
        when x"173A" => data_out<= x"00";
        when x"173B" => data_out<= x"20";
        when x"173C" => data_out<= x"AD";
        when x"173D" => data_out<= x"B0";
        when x"173E" => data_out<= x"20";
        when x"173F" => data_out<= x"4D";
        when x"1740" => data_out<= x"AF";
        when x"1741" => data_out<= x"20";
        when x"1742" => data_out<= x"E2";
        when x"1743" => data_out<= x"AE";
        when x"1744" => data_out<= x"4C";
        when x"1745" => data_out<= x"F5";
        when x"1746" => data_out<= x"96";
        when x"1747" => data_out<= x"A9";
        when x"1748" => data_out<= x"02";
        when x"1749" => data_out<= x"20";
        when x"174A" => data_out<= x"69";
        when x"174B" => data_out<= x"AF";
        when x"174C" => data_out<= x"20";
        when x"174D" => data_out<= x"7B";
        when x"174E" => data_out<= x"B0";
        when x"174F" => data_out<= x"A0";
        when x"1750" => data_out<= x"45";
        when x"1751" => data_out<= x"20";
        when x"1752" => data_out<= x"4F";
        when x"1753" => data_out<= x"AF";
        when x"1754" => data_out<= x"20";
        when x"1755" => data_out<= x"3B";
        when x"1756" => data_out<= x"A8";
        when x"1757" => data_out<= x"A0";
        when x"1758" => data_out<= x"43";
        when x"1759" => data_out<= x"20";
        when x"175A" => data_out<= x"4F";
        when x"175B" => data_out<= x"AF";
        when x"175C" => data_out<= x"A0";
        when x"175D" => data_out<= x"44";
        when x"175E" => data_out<= x"20";
        when x"175F" => data_out<= x"04";
        when x"1760" => data_out<= x"AE";
        when x"1761" => data_out<= x"A0";
        when x"1762" => data_out<= x"45";
        when x"1763" => data_out<= x"20";
        when x"1764" => data_out<= x"4F";
        when x"1765" => data_out<= x"AF";
        when x"1766" => data_out<= x"A8";
        when x"1767" => data_out<= x"8A";
        when x"1768" => data_out<= x"29";
        when x"1769" => data_out<= x"03";
        when x"176A" => data_out<= x"AA";
        when x"176B" => data_out<= x"98";
        when x"176C" => data_out<= x"E0";
        when x"176D" => data_out<= x"00";
        when x"176E" => data_out<= x"D0";
        when x"176F" => data_out<= x"09";
        when x"1770" => data_out<= x"C9";
        when x"1771" => data_out<= x"00";
        when x"1772" => data_out<= x"D0";
        when x"1773" => data_out<= x"05";
        when x"1774" => data_out<= x"A9";
        when x"1775" => data_out<= x"2E";
        when x"1776" => data_out<= x"20";
        when x"1777" => data_out<= x"F0";
        when x"1778" => data_out<= x"80";
        when x"1779" => data_out<= x"A0";
        when x"177A" => data_out<= x"45";
        when x"177B" => data_out<= x"20";
        when x"177C" => data_out<= x"4F";
        when x"177D" => data_out<= x"AF";
        when x"177E" => data_out<= x"A0";
        when x"177F" => data_out<= x"47";
        when x"1780" => data_out<= x"D1";
        when x"1781" => data_out<= x"0C";
        when x"1782" => data_out<= x"8A";
        when x"1783" => data_out<= x"C8";
        when x"1784" => data_out<= x"F1";
        when x"1785" => data_out<= x"0C";
        when x"1786" => data_out<= x"B0";
        when x"1787" => data_out<= x"03";
        when x"1788" => data_out<= x"4C";
        when x"1789" => data_out<= x"CF";
        when x"178A" => data_out<= x"96";
        when x"178B" => data_out<= x"20";
        when x"178C" => data_out<= x"B9";
        when x"178D" => data_out<= x"A9";
        when x"178E" => data_out<= x"20";
        when x"178F" => data_out<= x"45";
        when x"1790" => data_out<= x"8C";
        when x"1791" => data_out<= x"A9";
        when x"1792" => data_out<= x"A4";
        when x"1793" => data_out<= x"A2";
        when x"1794" => data_out<= x"BC";
        when x"1795" => data_out<= x"20";
        when x"1796" => data_out<= x"22";
        when x"1797" => data_out<= x"81";
        when x"1798" => data_out<= x"A0";
        when x"1799" => data_out<= x"45";
        when x"179A" => data_out<= x"20";
        when x"179B" => data_out<= x"4F";
        when x"179C" => data_out<= x"AF";
        when x"179D" => data_out<= x"20";
        when x"179E" => data_out<= x"86";
        when x"179F" => data_out<= x"93";
        when x"17A0" => data_out<= x"A9";
        when x"17A1" => data_out<= x"34";
        when x"17A2" => data_out<= x"A2";
        when x"17A3" => data_out<= x"BC";
        when x"17A4" => data_out<= x"20";
        when x"17A5" => data_out<= x"22";
        when x"17A6" => data_out<= x"81";
        when x"17A7" => data_out<= x"20";
        when x"17A8" => data_out<= x"45";
        when x"17A9" => data_out<= x"8C";
        when x"17AA" => data_out<= x"A0";
        when x"17AB" => data_out<= x"4D";
        when x"17AC" => data_out<= x"4C";
        when x"17AD" => data_out<= x"14";
        when x"17AE" => data_out<= x"AE";
        when x"17AF" => data_out<= x"20";
        when x"17B0" => data_out<= x"7B";
        when x"17B1" => data_out<= x"B0";
        when x"17B2" => data_out<= x"20";
        when x"17B3" => data_out<= x"6A";
        when x"17B4" => data_out<= x"AE";
        when x"17B5" => data_out<= x"20";
        when x"17B6" => data_out<= x"77";
        when x"17B7" => data_out<= x"B0";
        when x"17B8" => data_out<= x"A0";
        when x"17B9" => data_out<= x"46";
        when x"17BA" => data_out<= x"20";
        when x"17BB" => data_out<= x"13";
        when x"17BC" => data_out<= x"B1";
        when x"17BD" => data_out<= x"AD";
        when x"17BE" => data_out<= x"03";
        when x"17BF" => data_out<= x"02";
        when x"17C0" => data_out<= x"D0";
        when x"17C1" => data_out<= x"0D";
        when x"17C2" => data_out<= x"A9";
        when x"17C3" => data_out<= x"46";
        when x"17C4" => data_out<= x"A2";
        when x"17C5" => data_out<= x"BB";
        when x"17C6" => data_out<= x"20";
        when x"17C7" => data_out<= x"22";
        when x"17C8" => data_out<= x"81";
        when x"17C9" => data_out<= x"20";
        when x"17CA" => data_out<= x"45";
        when x"17CB" => data_out<= x"8C";
        when x"17CC" => data_out<= x"4C";
        when x"17CD" => data_out<= x"25";
        when x"17CE" => data_out<= x"99";
        when x"17CF" => data_out<= x"A0";
        when x"17D0" => data_out<= x"4C";
        when x"17D1" => data_out<= x"20";
        when x"17D2" => data_out<= x"4F";
        when x"17D3" => data_out<= x"AF";
        when x"17D4" => data_out<= x"20";
        when x"17D5" => data_out<= x"E0";
        when x"17D6" => data_out<= x"A3";
        when x"17D7" => data_out<= x"A0";
        when x"17D8" => data_out<= x"48";
        when x"17D9" => data_out<= x"91";
        when x"17DA" => data_out<= x"0C";
        when x"17DB" => data_out<= x"B1";
        when x"17DC" => data_out<= x"0C";
        when x"17DD" => data_out<= x"F0";
        when x"17DE" => data_out<= x"15";
        when x"17DF" => data_out<= x"A9";
        when x"17E0" => data_out<= x"C7";
        when x"17E1" => data_out<= x"A2";
        when x"17E2" => data_out<= x"BA";
        when x"17E3" => data_out<= x"20";
        when x"17E4" => data_out<= x"22";
        when x"17E5" => data_out<= x"81";
        when x"17E6" => data_out<= x"A0";
        when x"17E7" => data_out<= x"4C";
        when x"17E8" => data_out<= x"20";
        when x"17E9" => data_out<= x"4F";
        when x"17EA" => data_out<= x"AF";
        when x"17EB" => data_out<= x"20";
        when x"17EC" => data_out<= x"22";
        when x"17ED" => data_out<= x"81";
        when x"17EE" => data_out<= x"20";
        when x"17EF" => data_out<= x"45";
        when x"17F0" => data_out<= x"8C";
        when x"17F1" => data_out<= x"4C";
        when x"17F2" => data_out<= x"25";
        when x"17F3" => data_out<= x"99";
        when x"17F4" => data_out<= x"20";
        when x"17F5" => data_out<= x"30";
        when x"17F6" => data_out<= x"AB";
        when x"17F7" => data_out<= x"20";
        when x"17F8" => data_out<= x"C3";
        when x"17F9" => data_out<= x"B0";
        when x"17FA" => data_out<= x"A9";
        when x"17FB" => data_out<= x"EC";
        when x"17FC" => data_out<= x"A2";
        when x"17FD" => data_out<= x"BB";
        when x"17FE" => data_out<= x"20";
        when x"17FF" => data_out<= x"22";
        when x"1800" => data_out<= x"81";
        when x"1801" => data_out<= x"A0";
        when x"1802" => data_out<= x"4C";
        when x"1803" => data_out<= x"20";
        when x"1804" => data_out<= x"4F";
        when x"1805" => data_out<= x"AF";
        when x"1806" => data_out<= x"20";
        when x"1807" => data_out<= x"22";
        when x"1808" => data_out<= x"81";
        when x"1809" => data_out<= x"A9";
        when x"180A" => data_out<= x"F7";
        when x"180B" => data_out<= x"A2";
        when x"180C" => data_out<= x"B6";
        when x"180D" => data_out<= x"20";
        when x"180E" => data_out<= x"22";
        when x"180F" => data_out<= x"81";
        when x"1810" => data_out<= x"20";
        when x"1811" => data_out<= x"4D";
        when x"1812" => data_out<= x"AF";
        when x"1813" => data_out<= x"20";
        when x"1814" => data_out<= x"86";
        when x"1815" => data_out<= x"93";
        when x"1816" => data_out<= x"A9";
        when x"1817" => data_out<= x"8A";
        when x"1818" => data_out<= x"A2";
        when x"1819" => data_out<= x"BB";
        when x"181A" => data_out<= x"20";
        when x"181B" => data_out<= x"22";
        when x"181C" => data_out<= x"81";
        when x"181D" => data_out<= x"A0";
        when x"181E" => data_out<= x"4A";
        when x"181F" => data_out<= x"20";
        when x"1820" => data_out<= x"4F";
        when x"1821" => data_out<= x"AF";
        when x"1822" => data_out<= x"20";
        when x"1823" => data_out<= x"31";
        when x"1824" => data_out<= x"8C";
        when x"1825" => data_out<= x"20";
        when x"1826" => data_out<= x"45";
        when x"1827" => data_out<= x"8C";
        when x"1828" => data_out<= x"4C";
        when x"1829" => data_out<= x"C3";
        when x"182A" => data_out<= x"98";
        when x"182B" => data_out<= x"A9";
        when x"182C" => data_out<= x"04";
        when x"182D" => data_out<= x"20";
        when x"182E" => data_out<= x"69";
        when x"182F" => data_out<= x"AF";
        when x"1830" => data_out<= x"20";
        when x"1831" => data_out<= x"7B";
        when x"1832" => data_out<= x"B0";
        when x"1833" => data_out<= x"A2";
        when x"1834" => data_out<= x"00";
        when x"1835" => data_out<= x"A9";
        when x"1836" => data_out<= x"40";
        when x"1837" => data_out<= x"20";
        when x"1838" => data_out<= x"92";
        when x"1839" => data_out<= x"A6";
        when x"183A" => data_out<= x"A0";
        when x"183B" => data_out<= x"44";
        when x"183C" => data_out<= x"20";
        when x"183D" => data_out<= x"C5";
        when x"183E" => data_out<= x"B0";
        when x"183F" => data_out<= x"E0";
        when x"1840" => data_out<= x"00";
        when x"1841" => data_out<= x"D0";
        when x"1842" => data_out<= x"07";
        when x"1843" => data_out<= x"C9";
        when x"1844" => data_out<= x"00";
        when x"1845" => data_out<= x"D0";
        when x"1846" => data_out<= x"03";
        when x"1847" => data_out<= x"4C";
        when x"1848" => data_out<= x"D5";
        when x"1849" => data_out<= x"98";
        when x"184A" => data_out<= x"A2";
        when x"184B" => data_out<= x"00";
        when x"184C" => data_out<= x"8A";
        when x"184D" => data_out<= x"A0";
        when x"184E" => data_out<= x"02";
        when x"184F" => data_out<= x"20";
        when x"1850" => data_out<= x"C5";
        when x"1851" => data_out<= x"B0";
        when x"1852" => data_out<= x"A0";
        when x"1853" => data_out<= x"44";
        when x"1854" => data_out<= x"D1";
        when x"1855" => data_out<= x"0C";
        when x"1856" => data_out<= x"8A";
        when x"1857" => data_out<= x"C8";
        when x"1858" => data_out<= x"F1";
        when x"1859" => data_out<= x"0C";
        when x"185A" => data_out<= x"B0";
        when x"185B" => data_out<= x"47";
        when x"185C" => data_out<= x"A0";
        when x"185D" => data_out<= x"47";
        when x"185E" => data_out<= x"20";
        when x"185F" => data_out<= x"4F";
        when x"1860" => data_out<= x"AF";
        when x"1861" => data_out<= x"18";
        when x"1862" => data_out<= x"A0";
        when x"1863" => data_out<= x"49";
        when x"1864" => data_out<= x"71";
        when x"1865" => data_out<= x"0C";
        when x"1866" => data_out<= x"85";
        when x"1867" => data_out<= x"14";
        when x"1868" => data_out<= x"8A";
        when x"1869" => data_out<= x"C8";
        when x"186A" => data_out<= x"71";
        when x"186B" => data_out<= x"0C";
        when x"186C" => data_out<= x"85";
        when x"186D" => data_out<= x"15";
        when x"186E" => data_out<= x"A0";
        when x"186F" => data_out<= x"03";
        when x"1870" => data_out<= x"20";
        when x"1871" => data_out<= x"4F";
        when x"1872" => data_out<= x"AF";
        when x"1873" => data_out<= x"18";
        when x"1874" => data_out<= x"65";
        when x"1875" => data_out<= x"14";
        when x"1876" => data_out<= x"48";
        when x"1877" => data_out<= x"8A";
        when x"1878" => data_out<= x"65";
        when x"1879" => data_out<= x"15";
        when x"187A" => data_out<= x"AA";
        when x"187B" => data_out<= x"68";
        when x"187C" => data_out<= x"20";
        when x"187D" => data_out<= x"7B";
        when x"187E" => data_out<= x"B0";
        when x"187F" => data_out<= x"A9";
        when x"1880" => data_out<= x"06";
        when x"1881" => data_out<= x"20";
        when x"1882" => data_out<= x"69";
        when x"1883" => data_out<= x"AF";
        when x"1884" => data_out<= x"A0";
        when x"1885" => data_out<= x"04";
        when x"1886" => data_out<= x"18";
        when x"1887" => data_out<= x"71";
        when x"1888" => data_out<= x"0C";
        when x"1889" => data_out<= x"85";
        when x"188A" => data_out<= x"14";
        when x"188B" => data_out<= x"8A";
        when x"188C" => data_out<= x"C8";
        when x"188D" => data_out<= x"71";
        when x"188E" => data_out<= x"0C";
        when x"188F" => data_out<= x"85";
        when x"1890" => data_out<= x"15";
        when x"1891" => data_out<= x"A0";
        when x"1892" => data_out<= x"00";
        when x"1893" => data_out<= x"B1";
        when x"1894" => data_out<= x"14";
        when x"1895" => data_out<= x"20";
        when x"1896" => data_out<= x"5A";
        when x"1897" => data_out<= x"89";
        when x"1898" => data_out<= x"A0";
        when x"1899" => data_out<= x"03";
        when x"189A" => data_out<= x"20";
        when x"189B" => data_out<= x"4F";
        when x"189C" => data_out<= x"AF";
        when x"189D" => data_out<= x"20";
        when x"189E" => data_out<= x"E2";
        when x"189F" => data_out<= x"AE";
        when x"18A0" => data_out<= x"4C";
        when x"18A1" => data_out<= x"4D";
        when x"18A2" => data_out<= x"98";
        when x"18A3" => data_out<= x"20";
        when x"18A4" => data_out<= x"4F";
        when x"18A5" => data_out<= x"AF";
        when x"18A6" => data_out<= x"A0";
        when x"18A7" => data_out<= x"46";
        when x"18A8" => data_out<= x"20";
        when x"18A9" => data_out<= x"04";
        when x"18AA" => data_out<= x"AE";
        when x"18AB" => data_out<= x"A0";
        when x"18AC" => data_out<= x"47";
        when x"18AD" => data_out<= x"20";
        when x"18AE" => data_out<= x"4F";
        when x"18AF" => data_out<= x"AF";
        when x"18B0" => data_out<= x"A8";
        when x"18B1" => data_out<= x"8A";
        when x"18B2" => data_out<= x"29";
        when x"18B3" => data_out<= x"03";
        when x"18B4" => data_out<= x"AA";
        when x"18B5" => data_out<= x"98";
        when x"18B6" => data_out<= x"E0";
        when x"18B7" => data_out<= x"00";
        when x"18B8" => data_out<= x"D0";
        when x"18B9" => data_out<= x"09";
        when x"18BA" => data_out<= x"C9";
        when x"18BB" => data_out<= x"00";
        when x"18BC" => data_out<= x"D0";
        when x"18BD" => data_out<= x"05";
        when x"18BE" => data_out<= x"A9";
        when x"18BF" => data_out<= x"2E";
        when x"18C0" => data_out<= x"20";
        when x"18C1" => data_out<= x"F0";
        when x"18C2" => data_out<= x"80";
        when x"18C3" => data_out<= x"A0";
        when x"18C4" => data_out<= x"47";
        when x"18C5" => data_out<= x"20";
        when x"18C6" => data_out<= x"4F";
        when x"18C7" => data_out<= x"AF";
        when x"18C8" => data_out<= x"A0";
        when x"18C9" => data_out<= x"00";
        when x"18CA" => data_out<= x"D1";
        when x"18CB" => data_out<= x"0C";
        when x"18CC" => data_out<= x"8A";
        when x"18CD" => data_out<= x"C8";
        when x"18CE" => data_out<= x"F1";
        when x"18CF" => data_out<= x"0C";
        when x"18D0" => data_out<= x"B0";
        when x"18D1" => data_out<= x"03";
        when x"18D2" => data_out<= x"4C";
        when x"18D3" => data_out<= x"2B";
        when x"18D4" => data_out<= x"98";
        when x"18D5" => data_out<= x"20";
        when x"18D6" => data_out<= x"B9";
        when x"18D7" => data_out<= x"A9";
        when x"18D8" => data_out<= x"20";
        when x"18D9" => data_out<= x"45";
        when x"18DA" => data_out<= x"8C";
        when x"18DB" => data_out<= x"A9";
        when x"18DC" => data_out<= x"A4";
        when x"18DD" => data_out<= x"A2";
        when x"18DE" => data_out<= x"BC";
        when x"18DF" => data_out<= x"20";
        when x"18E0" => data_out<= x"22";
        when x"18E1" => data_out<= x"81";
        when x"18E2" => data_out<= x"A0";
        when x"18E3" => data_out<= x"47";
        when x"18E4" => data_out<= x"20";
        when x"18E5" => data_out<= x"4F";
        when x"18E6" => data_out<= x"AF";
        when x"18E7" => data_out<= x"20";
        when x"18E8" => data_out<= x"86";
        when x"18E9" => data_out<= x"93";
        when x"18EA" => data_out<= x"A9";
        when x"18EB" => data_out<= x"CA";
        when x"18EC" => data_out<= x"A2";
        when x"18ED" => data_out<= x"BB";
        when x"18EE" => data_out<= x"20";
        when x"18EF" => data_out<= x"22";
        when x"18F0" => data_out<= x"81";
        when x"18F1" => data_out<= x"A0";
        when x"18F2" => data_out<= x"4A";
        when x"18F3" => data_out<= x"20";
        when x"18F4" => data_out<= x"4F";
        when x"18F5" => data_out<= x"AF";
        when x"18F6" => data_out<= x"20";
        when x"18F7" => data_out<= x"31";
        when x"18F8" => data_out<= x"8C";
        when x"18F9" => data_out<= x"A9";
        when x"18FA" => data_out<= x"7D";
        when x"18FB" => data_out<= x"A2";
        when x"18FC" => data_out<= x"BD";
        when x"18FD" => data_out<= x"20";
        when x"18FE" => data_out<= x"22";
        when x"18FF" => data_out<= x"81";
        when x"1900" => data_out<= x"A0";
        when x"1901" => data_out<= x"47";
        when x"1902" => data_out<= x"20";
        when x"1903" => data_out<= x"4F";
        when x"1904" => data_out<= x"AF";
        when x"1905" => data_out<= x"18";
        when x"1906" => data_out<= x"A0";
        when x"1907" => data_out<= x"49";
        when x"1908" => data_out<= x"71";
        when x"1909" => data_out<= x"0C";
        when x"190A" => data_out<= x"48";
        when x"190B" => data_out<= x"8A";
        when x"190C" => data_out<= x"C8";
        when x"190D" => data_out<= x"71";
        when x"190E" => data_out<= x"0C";
        when x"190F" => data_out<= x"AA";
        when x"1910" => data_out<= x"68";
        when x"1911" => data_out<= x"20";
        when x"1912" => data_out<= x"5A";
        when x"1913" => data_out<= x"AE";
        when x"1914" => data_out<= x"20";
        when x"1915" => data_out<= x"31";
        when x"1916" => data_out<= x"8C";
        when x"1917" => data_out<= x"20";
        when x"1918" => data_out<= x"45";
        when x"1919" => data_out<= x"8C";
        when x"191A" => data_out<= x"A0";
        when x"191B" => data_out<= x"4A";
        when x"191C" => data_out<= x"20";
        when x"191D" => data_out<= x"4F";
        when x"191E" => data_out<= x"AF";
        when x"191F" => data_out<= x"8D";
        when x"1920" => data_out<= x"00";
        when x"1921" => data_out<= x"02";
        when x"1922" => data_out<= x"8E";
        when x"1923" => data_out<= x"01";
        when x"1924" => data_out<= x"02";
        when x"1925" => data_out<= x"A0";
        when x"1926" => data_out<= x"4D";
        when x"1927" => data_out<= x"4C";
        when x"1928" => data_out<= x"14";
        when x"1929" => data_out<= x"AE";
        when x"192A" => data_out<= x"20";
        when x"192B" => data_out<= x"7B";
        when x"192C" => data_out<= x"B0";
        when x"192D" => data_out<= x"20";
        when x"192E" => data_out<= x"6A";
        when x"192F" => data_out<= x"AE";
        when x"1930" => data_out<= x"AD";
        when x"1931" => data_out<= x"03";
        when x"1932" => data_out<= x"02";
        when x"1933" => data_out<= x"D0";
        when x"1934" => data_out<= x"0A";
        when x"1935" => data_out<= x"A9";
        when x"1936" => data_out<= x"46";
        when x"1937" => data_out<= x"A2";
        when x"1938" => data_out<= x"BB";
        when x"1939" => data_out<= x"20";
        when x"193A" => data_out<= x"22";
        when x"193B" => data_out<= x"81";
        when x"193C" => data_out<= x"4C";
        when x"193D" => data_out<= x"6F";
        when x"193E" => data_out<= x"99";
        when x"193F" => data_out<= x"A0";
        when x"1940" => data_out<= x"02";
        when x"1941" => data_out<= x"20";
        when x"1942" => data_out<= x"4F";
        when x"1943" => data_out<= x"AF";
        when x"1944" => data_out<= x"20";
        when x"1945" => data_out<= x"DF";
        when x"1946" => data_out<= x"A9";
        when x"1947" => data_out<= x"A0";
        when x"1948" => data_out<= x"00";
        when x"1949" => data_out<= x"91";
        when x"194A" => data_out<= x"0C";
        when x"194B" => data_out<= x"B1";
        when x"194C" => data_out<= x"0C";
        when x"194D" => data_out<= x"D0";
        when x"194E" => data_out<= x"12";
        when x"194F" => data_out<= x"A9";
        when x"1950" => data_out<= x"D6";
        when x"1951" => data_out<= x"A2";
        when x"1952" => data_out<= x"BB";
        when x"1953" => data_out<= x"20";
        when x"1954" => data_out<= x"22";
        when x"1955" => data_out<= x"81";
        when x"1956" => data_out<= x"A0";
        when x"1957" => data_out<= x"02";
        when x"1958" => data_out<= x"20";
        when x"1959" => data_out<= x"4F";
        when x"195A" => data_out<= x"AF";
        when x"195B" => data_out<= x"20";
        when x"195C" => data_out<= x"22";
        when x"195D" => data_out<= x"81";
        when x"195E" => data_out<= x"4C";
        when x"195F" => data_out<= x"6F";
        when x"1960" => data_out<= x"99";
        when x"1961" => data_out<= x"A9";
        when x"1962" => data_out<= x"2C";
        when x"1963" => data_out<= x"A2";
        when x"1964" => data_out<= x"BC";
        when x"1965" => data_out<= x"20";
        when x"1966" => data_out<= x"22";
        when x"1967" => data_out<= x"81";
        when x"1968" => data_out<= x"A0";
        when x"1969" => data_out<= x"00";
        when x"196A" => data_out<= x"B1";
        when x"196B" => data_out<= x"0C";
        when x"196C" => data_out<= x"20";
        when x"196D" => data_out<= x"FD";
        when x"196E" => data_out<= x"8B";
        when x"196F" => data_out<= x"20";
        when x"1970" => data_out<= x"45";
        when x"1971" => data_out<= x"8C";
        when x"1972" => data_out<= x"4C";
        when x"1973" => data_out<= x"22";
        when x"1974" => data_out<= x"AF";
        when x"1975" => data_out<= x"20";
        when x"1976" => data_out<= x"7B";
        when x"1977" => data_out<= x"B0";
        when x"1978" => data_out<= x"A0";
        when x"1979" => data_out<= x"11";
        when x"197A" => data_out<= x"20";
        when x"197B" => data_out<= x"13";
        when x"197C" => data_out<= x"B1";
        when x"197D" => data_out<= x"20";
        when x"197E" => data_out<= x"77";
        when x"197F" => data_out<= x"B0";
        when x"1980" => data_out<= x"20";
        when x"1981" => data_out<= x"80";
        when x"1982" => data_out<= x"AE";
        when x"1983" => data_out<= x"AD";
        when x"1984" => data_out<= x"03";
        when x"1985" => data_out<= x"02";
        when x"1986" => data_out<= x"D0";
        when x"1987" => data_out<= x"0D";
        when x"1988" => data_out<= x"A9";
        when x"1989" => data_out<= x"46";
        when x"198A" => data_out<= x"A2";
        when x"198B" => data_out<= x"BB";
        when x"198C" => data_out<= x"20";
        when x"198D" => data_out<= x"22";
        when x"198E" => data_out<= x"81";
        when x"198F" => data_out<= x"20";
        when x"1990" => data_out<= x"45";
        when x"1991" => data_out<= x"8C";
        when x"1992" => data_out<= x"4C";
        when x"1993" => data_out<= x"F4";
        when x"1994" => data_out<= x"9A";
        when x"1995" => data_out<= x"A0";
        when x"1996" => data_out<= x"17";
        when x"1997" => data_out<= x"20";
        when x"1998" => data_out<= x"4F";
        when x"1999" => data_out<= x"AF";
        when x"199A" => data_out<= x"20";
        when x"199B" => data_out<= x"E0";
        when x"199C" => data_out<= x"A3";
        when x"199D" => data_out<= x"A0";
        when x"199E" => data_out<= x"15";
        when x"199F" => data_out<= x"91";
        when x"19A0" => data_out<= x"0C";
        when x"19A1" => data_out<= x"B1";
        when x"19A2" => data_out<= x"0C";
        when x"19A3" => data_out<= x"F0";
        when x"19A4" => data_out<= x"0D";
        when x"19A5" => data_out<= x"A9";
        when x"19A6" => data_out<= x"54";
        when x"19A7" => data_out<= x"A2";
        when x"19A8" => data_out<= x"BB";
        when x"19A9" => data_out<= x"20";
        when x"19AA" => data_out<= x"22";
        when x"19AB" => data_out<= x"81";
        when x"19AC" => data_out<= x"20";
        when x"19AD" => data_out<= x"45";
        when x"19AE" => data_out<= x"8C";
        when x"19AF" => data_out<= x"4C";
        when x"19B0" => data_out<= x"F4";
        when x"19B1" => data_out<= x"9A";
        when x"19B2" => data_out<= x"A9";
        when x"19B3" => data_out<= x"B8";
        when x"19B4" => data_out<= x"A2";
        when x"19B5" => data_out<= x"BC";
        when x"19B6" => data_out<= x"20";
        when x"19B7" => data_out<= x"22";
        when x"19B8" => data_out<= x"81";
        when x"19B9" => data_out<= x"A0";
        when x"19BA" => data_out<= x"17";
        when x"19BB" => data_out<= x"20";
        when x"19BC" => data_out<= x"4F";
        when x"19BD" => data_out<= x"AF";
        when x"19BE" => data_out<= x"20";
        when x"19BF" => data_out<= x"22";
        when x"19C0" => data_out<= x"81";
        when x"19C1" => data_out<= x"A9";
        when x"19C2" => data_out<= x"B1";
        when x"19C3" => data_out<= x"A2";
        when x"19C4" => data_out<= x"B8";
        when x"19C5" => data_out<= x"20";
        when x"19C6" => data_out<= x"22";
        when x"19C7" => data_out<= x"81";
        when x"19C8" => data_out<= x"20";
        when x"19C9" => data_out<= x"45";
        when x"19CA" => data_out<= x"8C";
        when x"19CB" => data_out<= x"A9";
        when x"19CC" => data_out<= x"05";
        when x"19CD" => data_out<= x"20";
        when x"19CE" => data_out<= x"69";
        when x"19CF" => data_out<= x"AF";
        when x"19D0" => data_out<= x"20";
        when x"19D1" => data_out<= x"7B";
        when x"19D2" => data_out<= x"B0";
        when x"19D3" => data_out<= x"A2";
        when x"19D4" => data_out<= x"00";
        when x"19D5" => data_out<= x"A9";
        when x"19D6" => data_out<= x"10";
        when x"19D7" => data_out<= x"20";
        when x"19D8" => data_out<= x"92";
        when x"19D9" => data_out<= x"A6";
        when x"19DA" => data_out<= x"A0";
        when x"19DB" => data_out<= x"01";
        when x"19DC" => data_out<= x"20";
        when x"19DD" => data_out<= x"C5";
        when x"19DE" => data_out<= x"B0";
        when x"19DF" => data_out<= x"E0";
        when x"19E0" => data_out<= x"00";
        when x"19E1" => data_out<= x"D0";
        when x"19E2" => data_out<= x"07";
        when x"19E3" => data_out<= x"C9";
        when x"19E4" => data_out<= x"00";
        when x"19E5" => data_out<= x"D0";
        when x"19E6" => data_out<= x"03";
        when x"19E7" => data_out<= x"4C";
        when x"19E8" => data_out<= x"F1";
        when x"19E9" => data_out<= x"9A";
        when x"19EA" => data_out<= x"A0";
        when x"19EB" => data_out<= x"04";
        when x"19EC" => data_out<= x"20";
        when x"19ED" => data_out<= x"4F";
        when x"19EE" => data_out<= x"AF";
        when x"19EF" => data_out<= x"20";
        when x"19F0" => data_out<= x"31";
        when x"19F1" => data_out<= x"8C";
        when x"19F2" => data_out<= x"A9";
        when x"19F3" => data_out<= x"99";
        when x"19F4" => data_out<= x"A2";
        when x"19F5" => data_out<= x"B5";
        when x"19F6" => data_out<= x"20";
        when x"19F7" => data_out<= x"22";
        when x"19F8" => data_out<= x"81";
        when x"19F9" => data_out<= x"A9";
        when x"19FA" => data_out<= x"00";
        when x"19FB" => data_out<= x"A8";
        when x"19FC" => data_out<= x"91";
        when x"19FD" => data_out<= x"0C";
        when x"19FE" => data_out<= x"AA";
        when x"19FF" => data_out<= x"B1";
        when x"1A00" => data_out<= x"0C";
        when x"1A01" => data_out<= x"C8";
        when x"1A02" => data_out<= x"D1";
        when x"1A03" => data_out<= x"0C";
        when x"1A04" => data_out<= x"8A";
        when x"1A05" => data_out<= x"C8";
        when x"1A06" => data_out<= x"F1";
        when x"1A07" => data_out<= x"0C";
        when x"1A08" => data_out<= x"B0";
        when x"1A09" => data_out<= x"29";
        when x"1A0A" => data_out<= x"A9";
        when x"1A0B" => data_out<= x"05";
        when x"1A0C" => data_out<= x"20";
        when x"1A0D" => data_out<= x"69";
        when x"1A0E" => data_out<= x"AF";
        when x"1A0F" => data_out<= x"A0";
        when x"1A10" => data_out<= x"00";
        when x"1A11" => data_out<= x"18";
        when x"1A12" => data_out<= x"71";
        when x"1A13" => data_out<= x"0C";
        when x"1A14" => data_out<= x"90";
        when x"1A15" => data_out<= x"01";
        when x"1A16" => data_out<= x"E8";
        when x"1A17" => data_out<= x"85";
        when x"1A18" => data_out<= x"14";
        when x"1A19" => data_out<= x"86";
        when x"1A1A" => data_out<= x"15";
        when x"1A1B" => data_out<= x"B1";
        when x"1A1C" => data_out<= x"14";
        when x"1A1D" => data_out<= x"20";
        when x"1A1E" => data_out<= x"FD";
        when x"1A1F" => data_out<= x"8B";
        when x"1A20" => data_out<= x"A9";
        when x"1A21" => data_out<= x"20";
        when x"1A22" => data_out<= x"20";
        when x"1A23" => data_out<= x"F0";
        when x"1A24" => data_out<= x"80";
        when x"1A25" => data_out<= x"A0";
        when x"1A26" => data_out<= x"00";
        when x"1A27" => data_out<= x"A2";
        when x"1A28" => data_out<= x"00";
        when x"1A29" => data_out<= x"B1";
        when x"1A2A" => data_out<= x"0C";
        when x"1A2B" => data_out<= x"18";
        when x"1A2C" => data_out<= x"69";
        when x"1A2D" => data_out<= x"01";
        when x"1A2E" => data_out<= x"91";
        when x"1A2F" => data_out<= x"0C";
        when x"1A30" => data_out<= x"4C";
        when x"1A31" => data_out<= x"FF";
        when x"1A32" => data_out<= x"99";
        when x"1A33" => data_out<= x"A0";
        when x"1A34" => data_out<= x"00";
        when x"1A35" => data_out<= x"B1";
        when x"1A36" => data_out<= x"0C";
        when x"1A37" => data_out<= x"C9";
        when x"1A38" => data_out<= x"10";
        when x"1A39" => data_out<= x"B0";
        when x"1A3A" => data_out<= x"13";
        when x"1A3B" => data_out<= x"A9";
        when x"1A3C" => data_out<= x"01";
        when x"1A3D" => data_out<= x"A2";
        when x"1A3E" => data_out<= x"BD";
        when x"1A3F" => data_out<= x"20";
        when x"1A40" => data_out<= x"22";
        when x"1A41" => data_out<= x"81";
        when x"1A42" => data_out<= x"A0";
        when x"1A43" => data_out<= x"00";
        when x"1A44" => data_out<= x"B1";
        when x"1A45" => data_out<= x"0C";
        when x"1A46" => data_out<= x"18";
        when x"1A47" => data_out<= x"69";
        when x"1A48" => data_out<= x"01";
        when x"1A49" => data_out<= x"91";
        when x"1A4A" => data_out<= x"0C";
        when x"1A4B" => data_out<= x"4C";
        when x"1A4C" => data_out<= x"35";
        when x"1A4D" => data_out<= x"9A";
        when x"1A4E" => data_out<= x"A9";
        when x"1A4F" => data_out<= x"7C";
        when x"1A50" => data_out<= x"20";
        when x"1A51" => data_out<= x"F0";
        when x"1A52" => data_out<= x"80";
        when x"1A53" => data_out<= x"A9";
        when x"1A54" => data_out<= x"00";
        when x"1A55" => data_out<= x"A8";
        when x"1A56" => data_out<= x"91";
        when x"1A57" => data_out<= x"0C";
        when x"1A58" => data_out<= x"AA";
        when x"1A59" => data_out<= x"B1";
        when x"1A5A" => data_out<= x"0C";
        when x"1A5B" => data_out<= x"C8";
        when x"1A5C" => data_out<= x"D1";
        when x"1A5D" => data_out<= x"0C";
        when x"1A5E" => data_out<= x"8A";
        when x"1A5F" => data_out<= x"C8";
        when x"1A60" => data_out<= x"F1";
        when x"1A61" => data_out<= x"0C";
        when x"1A62" => data_out<= x"B0";
        when x"1A63" => data_out<= x"53";
        when x"1A64" => data_out<= x"A9";
        when x"1A65" => data_out<= x"05";
        when x"1A66" => data_out<= x"20";
        when x"1A67" => data_out<= x"69";
        when x"1A68" => data_out<= x"AF";
        when x"1A69" => data_out<= x"A0";
        when x"1A6A" => data_out<= x"00";
        when x"1A6B" => data_out<= x"18";
        when x"1A6C" => data_out<= x"71";
        when x"1A6D" => data_out<= x"0C";
        when x"1A6E" => data_out<= x"90";
        when x"1A6F" => data_out<= x"01";
        when x"1A70" => data_out<= x"E8";
        when x"1A71" => data_out<= x"85";
        when x"1A72" => data_out<= x"14";
        when x"1A73" => data_out<= x"86";
        when x"1A74" => data_out<= x"15";
        when x"1A75" => data_out<= x"B1";
        when x"1A76" => data_out<= x"14";
        when x"1A77" => data_out<= x"C9";
        when x"1A78" => data_out<= x"20";
        when x"1A79" => data_out<= x"90";
        when x"1A7A" => data_out<= x"29";
        when x"1A7B" => data_out<= x"A9";
        when x"1A7C" => data_out<= x"05";
        when x"1A7D" => data_out<= x"20";
        when x"1A7E" => data_out<= x"69";
        when x"1A7F" => data_out<= x"AF";
        when x"1A80" => data_out<= x"18";
        when x"1A81" => data_out<= x"71";
        when x"1A82" => data_out<= x"0C";
        when x"1A83" => data_out<= x"90";
        when x"1A84" => data_out<= x"01";
        when x"1A85" => data_out<= x"E8";
        when x"1A86" => data_out<= x"85";
        when x"1A87" => data_out<= x"14";
        when x"1A88" => data_out<= x"86";
        when x"1A89" => data_out<= x"15";
        when x"1A8A" => data_out<= x"B1";
        when x"1A8B" => data_out<= x"14";
        when x"1A8C" => data_out<= x"C9";
        when x"1A8D" => data_out<= x"7F";
        when x"1A8E" => data_out<= x"B0";
        when x"1A8F" => data_out<= x"14";
        when x"1A90" => data_out<= x"A9";
        when x"1A91" => data_out<= x"05";
        when x"1A92" => data_out<= x"20";
        when x"1A93" => data_out<= x"69";
        when x"1A94" => data_out<= x"AF";
        when x"1A95" => data_out<= x"18";
        when x"1A96" => data_out<= x"71";
        when x"1A97" => data_out<= x"0C";
        when x"1A98" => data_out<= x"90";
        when x"1A99" => data_out<= x"01";
        when x"1A9A" => data_out<= x"E8";
        when x"1A9B" => data_out<= x"85";
        when x"1A9C" => data_out<= x"14";
        when x"1A9D" => data_out<= x"86";
        when x"1A9E" => data_out<= x"15";
        when x"1A9F" => data_out<= x"B1";
        when x"1AA0" => data_out<= x"14";
        when x"1AA1" => data_out<= x"4C";
        when x"1AA2" => data_out<= x"A6";
        when x"1AA3" => data_out<= x"9A";
        when x"1AA4" => data_out<= x"A9";
        when x"1AA5" => data_out<= x"2E";
        when x"1AA6" => data_out<= x"20";
        when x"1AA7" => data_out<= x"F0";
        when x"1AA8" => data_out<= x"80";
        when x"1AA9" => data_out<= x"A0";
        when x"1AAA" => data_out<= x"00";
        when x"1AAB" => data_out<= x"A2";
        when x"1AAC" => data_out<= x"00";
        when x"1AAD" => data_out<= x"B1";
        when x"1AAE" => data_out<= x"0C";
        when x"1AAF" => data_out<= x"18";
        when x"1AB0" => data_out<= x"69";
        when x"1AB1" => data_out<= x"01";
        when x"1AB2" => data_out<= x"91";
        when x"1AB3" => data_out<= x"0C";
        when x"1AB4" => data_out<= x"4C";
        when x"1AB5" => data_out<= x"59";
        when x"1AB6" => data_out<= x"9A";
        when x"1AB7" => data_out<= x"A9";
        when x"1AB8" => data_out<= x"7C";
        when x"1AB9" => data_out<= x"20";
        when x"1ABA" => data_out<= x"F0";
        when x"1ABB" => data_out<= x"80";
        when x"1ABC" => data_out<= x"20";
        when x"1ABD" => data_out<= x"45";
        when x"1ABE" => data_out<= x"8C";
        when x"1ABF" => data_out<= x"A0";
        when x"1AC0" => data_out<= x"02";
        when x"1AC1" => data_out<= x"20";
        when x"1AC2" => data_out<= x"4F";
        when x"1AC3" => data_out<= x"AF";
        when x"1AC4" => data_out<= x"A0";
        when x"1AC5" => data_out<= x"03";
        when x"1AC6" => data_out<= x"20";
        when x"1AC7" => data_out<= x"04";
        when x"1AC8" => data_out<= x"AE";
        when x"1AC9" => data_out<= x"A0";
        when x"1ACA" => data_out<= x"04";
        when x"1ACB" => data_out<= x"20";
        when x"1ACC" => data_out<= x"4F";
        when x"1ACD" => data_out<= x"AF";
        when x"1ACE" => data_out<= x"C9";
        when x"1ACF" => data_out<= x"00";
        when x"1AD0" => data_out<= x"8A";
        when x"1AD1" => data_out<= x"E9";
        when x"1AD2" => data_out<= x"01";
        when x"1AD3" => data_out<= x"B0";
        when x"1AD4" => data_out<= x"03";
        when x"1AD5" => data_out<= x"4C";
        when x"1AD6" => data_out<= x"CB";
        when x"1AD7" => data_out<= x"99";
        when x"1AD8" => data_out<= x"A9";
        when x"1AD9" => data_out<= x"C7";
        when x"1ADA" => data_out<= x"A2";
        when x"1ADB" => data_out<= x"BC";
        when x"1ADC" => data_out<= x"20";
        when x"1ADD" => data_out<= x"22";
        when x"1ADE" => data_out<= x"81";
        when x"1ADF" => data_out<= x"A0";
        when x"1AE0" => data_out<= x"04";
        when x"1AE1" => data_out<= x"20";
        when x"1AE2" => data_out<= x"4F";
        when x"1AE3" => data_out<= x"AF";
        when x"1AE4" => data_out<= x"20";
        when x"1AE5" => data_out<= x"86";
        when x"1AE6" => data_out<= x"93";
        when x"1AE7" => data_out<= x"A9";
        when x"1AE8" => data_out<= x"70";
        when x"1AE9" => data_out<= x"A2";
        when x"1AEA" => data_out<= x"BA";
        when x"1AEB" => data_out<= x"20";
        when x"1AEC" => data_out<= x"22";
        when x"1AED" => data_out<= x"81";
        when x"1AEE" => data_out<= x"20";
        when x"1AEF" => data_out<= x"45";
        when x"1AF0" => data_out<= x"8C";
        when x"1AF1" => data_out<= x"20";
        when x"1AF2" => data_out<= x"B9";
        when x"1AF3" => data_out<= x"A9";
        when x"1AF4" => data_out<= x"A0";
        when x"1AF5" => data_out<= x"18";
        when x"1AF6" => data_out<= x"4C";
        when x"1AF7" => data_out<= x"14";
        when x"1AF8" => data_out<= x"AE";
        when x"1AF9" => data_out<= x"20";
        when x"1AFA" => data_out<= x"7B";
        when x"1AFB" => data_out<= x"B0";
        when x"1AFC" => data_out<= x"4C";
        when x"1AFD" => data_out<= x"5F";
        when x"1AFE" => data_out<= x"9B";
        when x"1AFF" => data_out<= x"A0";
        when x"1B00" => data_out<= x"03";
        when x"1B01" => data_out<= x"20";
        when x"1B02" => data_out<= x"4F";
        when x"1B03" => data_out<= x"AF";
        when x"1B04" => data_out<= x"85";
        when x"1B05" => data_out<= x"14";
        when x"1B06" => data_out<= x"86";
        when x"1B07" => data_out<= x"15";
        when x"1B08" => data_out<= x"A0";
        when x"1B09" => data_out<= x"00";
        when x"1B0A" => data_out<= x"B1";
        when x"1B0B" => data_out<= x"14";
        when x"1B0C" => data_out<= x"20";
        when x"1B0D" => data_out<= x"65";
        when x"1B0E" => data_out<= x"B0";
        when x"1B0F" => data_out<= x"A0";
        when x"1B10" => data_out<= x"00";
        when x"1B11" => data_out<= x"B1";
        when x"1B12" => data_out<= x"0C";
        when x"1B13" => data_out<= x"C9";
        when x"1B14" => data_out<= x"61";
        when x"1B15" => data_out<= x"90";
        when x"1B16" => data_out<= x"0B";
        when x"1B17" => data_out<= x"B1";
        when x"1B18" => data_out<= x"0C";
        when x"1B19" => data_out<= x"C9";
        when x"1B1A" => data_out<= x"7B";
        when x"1B1B" => data_out<= x"B0";
        when x"1B1C" => data_out<= x"05";
        when x"1B1D" => data_out<= x"38";
        when x"1B1E" => data_out<= x"E9";
        when x"1B1F" => data_out<= x"20";
        when x"1B20" => data_out<= x"91";
        when x"1B21" => data_out<= x"0C";
        when x"1B22" => data_out<= x"B1";
        when x"1B23" => data_out<= x"0C";
        when x"1B24" => data_out<= x"20";
        when x"1B25" => data_out<= x"79";
        when x"1B26" => data_out<= x"B0";
        when x"1B27" => data_out<= x"A0";
        when x"1B28" => data_out<= x"04";
        when x"1B29" => data_out<= x"20";
        when x"1B2A" => data_out<= x"4F";
        when x"1B2B" => data_out<= x"AF";
        when x"1B2C" => data_out<= x"85";
        when x"1B2D" => data_out<= x"14";
        when x"1B2E" => data_out<= x"86";
        when x"1B2F" => data_out<= x"15";
        when x"1B30" => data_out<= x"A2";
        when x"1B31" => data_out<= x"00";
        when x"1B32" => data_out<= x"A1";
        when x"1B33" => data_out<= x"14";
        when x"1B34" => data_out<= x"20";
        when x"1B35" => data_out<= x"B4";
        when x"1B36" => data_out<= x"AE";
        when x"1B37" => data_out<= x"F0";
        when x"1B38" => data_out<= x"09";
        when x"1B39" => data_out<= x"A2";
        when x"1B3A" => data_out<= x"00";
        when x"1B3B" => data_out<= x"8A";
        when x"1B3C" => data_out<= x"20";
        when x"1B3D" => data_out<= x"05";
        when x"1B3E" => data_out<= x"AF";
        when x"1B3F" => data_out<= x"4C";
        when x"1B40" => data_out<= x"27";
        when x"1B41" => data_out<= x"AF";
        when x"1B42" => data_out<= x"A0";
        when x"1B43" => data_out<= x"04";
        when x"1B44" => data_out<= x"20";
        when x"1B45" => data_out<= x"4F";
        when x"1B46" => data_out<= x"AF";
        when x"1B47" => data_out<= x"20";
        when x"1B48" => data_out<= x"E2";
        when x"1B49" => data_out<= x"AE";
        when x"1B4A" => data_out<= x"A0";
        when x"1B4B" => data_out<= x"03";
        when x"1B4C" => data_out<= x"20";
        when x"1B4D" => data_out<= x"C5";
        when x"1B4E" => data_out<= x"B0";
        when x"1B4F" => data_out<= x"A0";
        when x"1B50" => data_out<= x"02";
        when x"1B51" => data_out<= x"20";
        when x"1B52" => data_out<= x"4F";
        when x"1B53" => data_out<= x"AF";
        when x"1B54" => data_out<= x"20";
        when x"1B55" => data_out<= x"E2";
        when x"1B56" => data_out<= x"AE";
        when x"1B57" => data_out<= x"A0";
        when x"1B58" => data_out<= x"01";
        when x"1B59" => data_out<= x"20";
        when x"1B5A" => data_out<= x"C5";
        when x"1B5B" => data_out<= x"B0";
        when x"1B5C" => data_out<= x"20";
        when x"1B5D" => data_out<= x"05";
        when x"1B5E" => data_out<= x"AF";
        when x"1B5F" => data_out<= x"20";
        when x"1B60" => data_out<= x"4D";
        when x"1B61" => data_out<= x"AF";
        when x"1B62" => data_out<= x"85";
        when x"1B63" => data_out<= x"14";
        when x"1B64" => data_out<= x"86";
        when x"1B65" => data_out<= x"15";
        when x"1B66" => data_out<= x"A0";
        when x"1B67" => data_out<= x"00";
        when x"1B68" => data_out<= x"B1";
        when x"1B69" => data_out<= x"14";
        when x"1B6A" => data_out<= x"D0";
        when x"1B6B" => data_out<= x"93";
        when x"1B6C" => data_out<= x"A0";
        when x"1B6D" => data_out<= x"03";
        when x"1B6E" => data_out<= x"20";
        when x"1B6F" => data_out<= x"4F";
        when x"1B70" => data_out<= x"AF";
        when x"1B71" => data_out<= x"85";
        when x"1B72" => data_out<= x"14";
        when x"1B73" => data_out<= x"86";
        when x"1B74" => data_out<= x"15";
        when x"1B75" => data_out<= x"A0";
        when x"1B76" => data_out<= x"00";
        when x"1B77" => data_out<= x"B1";
        when x"1B78" => data_out<= x"14";
        when x"1B79" => data_out<= x"C9";
        when x"1B7A" => data_out<= x"20";
        when x"1B7B" => data_out<= x"F0";
        when x"1B7C" => data_out<= x"15";
        when x"1B7D" => data_out<= x"A0";
        when x"1B7E" => data_out<= x"03";
        when x"1B7F" => data_out<= x"20";
        when x"1B80" => data_out<= x"4F";
        when x"1B81" => data_out<= x"AF";
        when x"1B82" => data_out<= x"85";
        when x"1B83" => data_out<= x"14";
        when x"1B84" => data_out<= x"86";
        when x"1B85" => data_out<= x"15";
        when x"1B86" => data_out<= x"A0";
        when x"1B87" => data_out<= x"00";
        when x"1B88" => data_out<= x"B1";
        when x"1B89" => data_out<= x"14";
        when x"1B8A" => data_out<= x"F0";
        when x"1B8B" => data_out<= x"06";
        when x"1B8C" => data_out<= x"A2";
        when x"1B8D" => data_out<= x"00";
        when x"1B8E" => data_out<= x"8A";
        when x"1B8F" => data_out<= x"4C";
        when x"1B90" => data_out<= x"27";
        when x"1B91" => data_out<= x"AF";
        when x"1B92" => data_out<= x"A9";
        when x"1B93" => data_out<= x"01";
        when x"1B94" => data_out<= x"A2";
        when x"1B95" => data_out<= x"00";
        when x"1B96" => data_out<= x"4C";
        when x"1B97" => data_out<= x"27";
        when x"1B98" => data_out<= x"AF";
        when x"1B99" => data_out<= x"20";
        when x"1B9A" => data_out<= x"45";
        when x"1B9B" => data_out<= x"8C";
        when x"1B9C" => data_out<= x"A9";
        when x"1B9D" => data_out<= x"B6";
        when x"1B9E" => data_out<= x"A2";
        when x"1B9F" => data_out<= x"B8";
        when x"1BA0" => data_out<= x"20";
        when x"1BA1" => data_out<= x"22";
        when x"1BA2" => data_out<= x"81";
        when x"1BA3" => data_out<= x"A9";
        when x"1BA4" => data_out<= x"5A";
        when x"1BA5" => data_out<= x"A2";
        when x"1BA6" => data_out<= x"B2";
        when x"1BA7" => data_out<= x"20";
        when x"1BA8" => data_out<= x"22";
        when x"1BA9" => data_out<= x"81";
        when x"1BAA" => data_out<= x"A9";
        when x"1BAB" => data_out<= x"CD";
        when x"1BAC" => data_out<= x"A2";
        when x"1BAD" => data_out<= x"B8";
        when x"1BAE" => data_out<= x"20";
        when x"1BAF" => data_out<= x"22";
        when x"1BB0" => data_out<= x"81";
        when x"1BB1" => data_out<= x"A9";
        when x"1BB2" => data_out<= x"29";
        when x"1BB3" => data_out<= x"A2";
        when x"1BB4" => data_out<= x"B9";
        when x"1BB5" => data_out<= x"20";
        when x"1BB6" => data_out<= x"22";
        when x"1BB7" => data_out<= x"81";
        when x"1BB8" => data_out<= x"A9";
        when x"1BB9" => data_out<= x"55";
        when x"1BBA" => data_out<= x"A2";
        when x"1BBB" => data_out<= x"B9";
        when x"1BBC" => data_out<= x"20";
        when x"1BBD" => data_out<= x"22";
        when x"1BBE" => data_out<= x"81";
        when x"1BBF" => data_out<= x"A9";
        when x"1BC0" => data_out<= x"55";
        when x"1BC1" => data_out<= x"A2";
        when x"1BC2" => data_out<= x"B4";
        when x"1BC3" => data_out<= x"20";
        when x"1BC4" => data_out<= x"22";
        when x"1BC5" => data_out<= x"81";
        when x"1BC6" => data_out<= x"A9";
        when x"1BC7" => data_out<= x"45";
        when x"1BC8" => data_out<= x"A2";
        when x"1BC9" => data_out<= x"B5";
        when x"1BCA" => data_out<= x"20";
        when x"1BCB" => data_out<= x"22";
        when x"1BCC" => data_out<= x"81";
        when x"1BCD" => data_out<= x"A9";
        when x"1BCE" => data_out<= x"82";
        when x"1BCF" => data_out<= x"A2";
        when x"1BD0" => data_out<= x"BA";
        when x"1BD1" => data_out<= x"20";
        when x"1BD2" => data_out<= x"22";
        when x"1BD3" => data_out<= x"81";
        when x"1BD4" => data_out<= x"A9";
        when x"1BD5" => data_out<= x"62";
        when x"1BD6" => data_out<= x"A2";
        when x"1BD7" => data_out<= x"B7";
        when x"1BD8" => data_out<= x"20";
        when x"1BD9" => data_out<= x"22";
        when x"1BDA" => data_out<= x"81";
        when x"1BDB" => data_out<= x"A9";
        when x"1BDC" => data_out<= x"0D";
        when x"1BDD" => data_out<= x"A2";
        when x"1BDE" => data_out<= x"B3";
        when x"1BDF" => data_out<= x"20";
        when x"1BE0" => data_out<= x"22";
        when x"1BE1" => data_out<= x"81";
        when x"1BE2" => data_out<= x"A9";
        when x"1BE3" => data_out<= x"78";
        when x"1BE4" => data_out<= x"A2";
        when x"1BE5" => data_out<= x"B6";
        when x"1BE6" => data_out<= x"20";
        when x"1BE7" => data_out<= x"22";
        when x"1BE8" => data_out<= x"81";
        when x"1BE9" => data_out<= x"A9";
        when x"1BEA" => data_out<= x"7D";
        when x"1BEB" => data_out<= x"A2";
        when x"1BEC" => data_out<= x"BB";
        when x"1BED" => data_out<= x"20";
        when x"1BEE" => data_out<= x"22";
        when x"1BEF" => data_out<= x"81";
        when x"1BF0" => data_out<= x"A9";
        when x"1BF1" => data_out<= x"C8";
        when x"1BF2" => data_out<= x"A2";
        when x"1BF3" => data_out<= x"B2";
        when x"1BF4" => data_out<= x"20";
        when x"1BF5" => data_out<= x"22";
        when x"1BF6" => data_out<= x"81";
        when x"1BF7" => data_out<= x"A9";
        when x"1BF8" => data_out<= x"24";
        when x"1BF9" => data_out<= x"A2";
        when x"1BFA" => data_out<= x"BA";
        when x"1BFB" => data_out<= x"20";
        when x"1BFC" => data_out<= x"22";
        when x"1BFD" => data_out<= x"81";
        when x"1BFE" => data_out<= x"A9";
        when x"1BFF" => data_out<= x"86";
        when x"1C00" => data_out<= x"A2";
        when x"1C01" => data_out<= x"B8";
        when x"1C02" => data_out<= x"4C";
        when x"1C03" => data_out<= x"22";
        when x"1C04" => data_out<= x"81";
        when x"1C05" => data_out<= x"20";
        when x"1C06" => data_out<= x"65";
        when x"1C07" => data_out<= x"B0";
        when x"1C08" => data_out<= x"A0";
        when x"1C09" => data_out<= x"00";
        when x"1C0A" => data_out<= x"B1";
        when x"1C0B" => data_out<= x"0C";
        when x"1C0C" => data_out<= x"C9";
        when x"1C0D" => data_out<= x"61";
        when x"1C0E" => data_out<= x"90";
        when x"1C0F" => data_out<= x"09";
        when x"1C10" => data_out<= x"C9";
        when x"1C11" => data_out<= x"7B";
        when x"1C12" => data_out<= x"B0";
        when x"1C13" => data_out<= x"05";
        when x"1C14" => data_out<= x"38";
        when x"1C15" => data_out<= x"E9";
        when x"1C16" => data_out<= x"20";
        when x"1C17" => data_out<= x"91";
        when x"1C18" => data_out<= x"0C";
        when x"1C19" => data_out<= x"20";
        when x"1C1A" => data_out<= x"45";
        when x"1C1B" => data_out<= x"8C";
        when x"1C1C" => data_out<= x"A0";
        when x"1C1D" => data_out<= x"00";
        when x"1C1E" => data_out<= x"B1";
        when x"1C1F" => data_out<= x"0C";
        when x"1C20" => data_out<= x"C9";
        when x"1C21" => data_out<= x"44";
        when x"1C22" => data_out<= x"F0";
        when x"1C23" => data_out<= x"5D";
        when x"1C24" => data_out<= x"C9";
        when x"1C25" => data_out<= x"46";
        when x"1C26" => data_out<= x"F0";
        when x"1C27" => data_out<= x"7C";
        when x"1C28" => data_out<= x"C9";
        when x"1C29" => data_out<= x"49";
        when x"1C2A" => data_out<= x"D0";
        when x"1C2B" => data_out<= x"03";
        when x"1C2C" => data_out<= x"4C";
        when x"1C2D" => data_out<= x"C7";
        when x"1C2E" => data_out<= x"9C";
        when x"1C2F" => data_out<= x"C9";
        when x"1C30" => data_out<= x"4C";
        when x"1C31" => data_out<= x"F0";
        when x"1C32" => data_out<= x"5C";
        when x"1C33" => data_out<= x"C9";
        when x"1C34" => data_out<= x"4D";
        when x"1C35" => data_out<= x"F0";
        when x"1C36" => data_out<= x"7B";
        when x"1C37" => data_out<= x"C9";
        when x"1C38" => data_out<= x"51";
        when x"1C39" => data_out<= x"D0";
        when x"1C3A" => data_out<= x"03";
        when x"1C3B" => data_out<= x"4C";
        when x"1C3C" => data_out<= x"D5";
        when x"1C3D" => data_out<= x"9C";
        when x"1C3E" => data_out<= x"C9";
        when x"1C3F" => data_out<= x"52";
        when x"1C40" => data_out<= x"F0";
        when x"1C41" => data_out<= x"07";
        when x"1C42" => data_out<= x"C9";
        when x"1C43" => data_out<= x"57";
        when x"1C44" => data_out<= x"F0";
        when x"1C45" => data_out<= x"2D";
        when x"1C46" => data_out<= x"4C";
        when x"1C47" => data_out<= x"DC";
        when x"1C48" => data_out<= x"9C";
        when x"1C49" => data_out<= x"A9";
        when x"1C4A" => data_out<= x"B4";
        when x"1C4B" => data_out<= x"A2";
        when x"1C4C" => data_out<= x"B3";
        when x"1C4D" => data_out<= x"20";
        when x"1C4E" => data_out<= x"22";
        when x"1C4F" => data_out<= x"81";
        when x"1C50" => data_out<= x"A9";
        when x"1C51" => data_out<= x"AB";
        when x"1C52" => data_out<= x"A2";
        when x"1C53" => data_out<= x"B9";
        when x"1C54" => data_out<= x"20";
        when x"1C55" => data_out<= x"22";
        when x"1C56" => data_out<= x"81";
        when x"1C57" => data_out<= x"A9";
        when x"1C58" => data_out<= x"93";
        when x"1C59" => data_out<= x"A2";
        when x"1C5A" => data_out<= x"B4";
        when x"1C5B" => data_out<= x"20";
        when x"1C5C" => data_out<= x"22";
        when x"1C5D" => data_out<= x"81";
        when x"1C5E" => data_out<= x"A9";
        when x"1C5F" => data_out<= x"26";
        when x"1C60" => data_out<= x"A2";
        when x"1C61" => data_out<= x"B8";
        when x"1C62" => data_out<= x"20";
        when x"1C63" => data_out<= x"22";
        when x"1C64" => data_out<= x"81";
        when x"1C65" => data_out<= x"A9";
        when x"1C66" => data_out<= x"6B";
        when x"1C67" => data_out<= x"A2";
        when x"1C68" => data_out<= x"B9";
        when x"1C69" => data_out<= x"20";
        when x"1C6A" => data_out<= x"22";
        when x"1C6B" => data_out<= x"81";
        when x"1C6C" => data_out<= x"A9";
        when x"1C6D" => data_out<= x"E4";
        when x"1C6E" => data_out<= x"A2";
        when x"1C6F" => data_out<= x"B8";
        when x"1C70" => data_out<= x"4C";
        when x"1C71" => data_out<= x"EE";
        when x"1C72" => data_out<= x"9C";
        when x"1C73" => data_out<= x"A9";
        when x"1C74" => data_out<= x"28";
        when x"1C75" => data_out<= x"A2";
        when x"1C76" => data_out<= x"B5";
        when x"1C77" => data_out<= x"20";
        when x"1C78" => data_out<= x"22";
        when x"1C79" => data_out<= x"81";
        when x"1C7A" => data_out<= x"A9";
        when x"1C7B" => data_out<= x"5D";
        when x"1C7C" => data_out<= x"A2";
        when x"1C7D" => data_out<= x"B6";
        when x"1C7E" => data_out<= x"4C";
        when x"1C7F" => data_out<= x"EE";
        when x"1C80" => data_out<= x"9C";
        when x"1C81" => data_out<= x"A9";
        when x"1C82" => data_out<= x"D5";
        when x"1C83" => data_out<= x"A2";
        when x"1C84" => data_out<= x"B3";
        when x"1C85" => data_out<= x"20";
        when x"1C86" => data_out<= x"22";
        when x"1C87" => data_out<= x"81";
        when x"1C88" => data_out<= x"A9";
        when x"1C89" => data_out<= x"51";
        when x"1C8A" => data_out<= x"A2";
        when x"1C8B" => data_out<= x"B3";
        when x"1C8C" => data_out<= x"4C";
        when x"1C8D" => data_out<= x"EE";
        when x"1C8E" => data_out<= x"9C";
        when x"1C8F" => data_out<= x"A9";
        when x"1C90" => data_out<= x"EB";
        when x"1C91" => data_out<= x"A2";
        when x"1C92" => data_out<= x"B2";
        when x"1C93" => data_out<= x"20";
        when x"1C94" => data_out<= x"22";
        when x"1C95" => data_out<= x"81";
        when x"1C96" => data_out<= x"A9";
        when x"1C97" => data_out<= x"9C";
        when x"1C98" => data_out<= x"A2";
        when x"1C99" => data_out<= x"B5";
        when x"1C9A" => data_out<= x"20";
        when x"1C9B" => data_out<= x"22";
        when x"1C9C" => data_out<= x"81";
        when x"1C9D" => data_out<= x"A9";
        when x"1C9E" => data_out<= x"A4";
        when x"1C9F" => data_out<= x"A2";
        when x"1CA0" => data_out<= x"B2";
        when x"1CA1" => data_out<= x"4C";
        when x"1CA2" => data_out<= x"EE";
        when x"1CA3" => data_out<= x"9C";
        when x"1CA4" => data_out<= x"A9";
        when x"1CA5" => data_out<= x"15";
        when x"1CA6" => data_out<= x"A2";
        when x"1CA7" => data_out<= x"B4";
        when x"1CA8" => data_out<= x"20";
        when x"1CA9" => data_out<= x"22";
        when x"1CAA" => data_out<= x"81";
        when x"1CAB" => data_out<= x"A9";
        when x"1CAC" => data_out<= x"2F";
        when x"1CAD" => data_out<= x"A2";
        when x"1CAE" => data_out<= x"B3";
        when x"1CAF" => data_out<= x"4C";
        when x"1CB0" => data_out<= x"EE";
        when x"1CB1" => data_out<= x"9C";
        when x"1CB2" => data_out<= x"A9";
        when x"1CB3" => data_out<= x"B9";
        when x"1CB4" => data_out<= x"A2";
        when x"1CB5" => data_out<= x"B5";
        when x"1CB6" => data_out<= x"20";
        when x"1CB7" => data_out<= x"22";
        when x"1CB8" => data_out<= x"81";
        when x"1CB9" => data_out<= x"A9";
        when x"1CBA" => data_out<= x"F1";
        when x"1CBB" => data_out<= x"A2";
        when x"1CBC" => data_out<= x"B5";
        when x"1CBD" => data_out<= x"20";
        when x"1CBE" => data_out<= x"22";
        when x"1CBF" => data_out<= x"81";
        when x"1CC0" => data_out<= x"A9";
        when x"1CC1" => data_out<= x"DE";
        when x"1CC2" => data_out<= x"A2";
        when x"1CC3" => data_out<= x"B7";
        when x"1CC4" => data_out<= x"4C";
        when x"1CC5" => data_out<= x"EE";
        when x"1CC6" => data_out<= x"9C";
        when x"1CC7" => data_out<= x"A9";
        when x"1CC8" => data_out<= x"F6";
        when x"1CC9" => data_out<= x"A2";
        when x"1CCA" => data_out<= x"B7";
        when x"1CCB" => data_out<= x"20";
        when x"1CCC" => data_out<= x"22";
        when x"1CCD" => data_out<= x"81";
        when x"1CCE" => data_out<= x"A9";
        when x"1CCF" => data_out<= x"0D";
        when x"1CD0" => data_out<= x"A2";
        when x"1CD1" => data_out<= x"B2";
        when x"1CD2" => data_out<= x"4C";
        when x"1CD3" => data_out<= x"EE";
        when x"1CD4" => data_out<= x"9C";
        when x"1CD5" => data_out<= x"A9";
        when x"1CD6" => data_out<= x"0E";
        when x"1CD7" => data_out<= x"A2";
        when x"1CD8" => data_out<= x"B8";
        when x"1CD9" => data_out<= x"4C";
        when x"1CDA" => data_out<= x"EE";
        when x"1CDB" => data_out<= x"9C";
        when x"1CDC" => data_out<= x"A9";
        when x"1CDD" => data_out<= x"49";
        when x"1CDE" => data_out<= x"A2";
        when x"1CDF" => data_out<= x"BC";
        when x"1CE0" => data_out<= x"20";
        when x"1CE1" => data_out<= x"22";
        when x"1CE2" => data_out<= x"81";
        when x"1CE3" => data_out<= x"A0";
        when x"1CE4" => data_out<= x"00";
        when x"1CE5" => data_out<= x"B1";
        when x"1CE6" => data_out<= x"0C";
        when x"1CE7" => data_out<= x"20";
        when x"1CE8" => data_out<= x"F0";
        when x"1CE9" => data_out<= x"80";
        when x"1CEA" => data_out<= x"A9";
        when x"1CEB" => data_out<= x"81";
        when x"1CEC" => data_out<= x"A2";
        when x"1CED" => data_out<= x"B9";
        when x"1CEE" => data_out<= x"20";
        when x"1CEF" => data_out<= x"22";
        when x"1CF0" => data_out<= x"81";
        when x"1CF1" => data_out<= x"4C";
        when x"1CF2" => data_out<= x"05";
        when x"1CF3" => data_out<= x"AF";
        when x"1CF4" => data_out<= x"20";
        when x"1CF5" => data_out<= x"7B";
        when x"1CF6" => data_out<= x"B0";
        when x"1CF7" => data_out<= x"20";
        when x"1CF8" => data_out<= x"45";
        when x"1CF9" => data_out<= x"8C";
        when x"1CFA" => data_out<= x"20";
        when x"1CFB" => data_out<= x"91";
        when x"1CFC" => data_out<= x"B0";
        when x"1CFD" => data_out<= x"A9";
        when x"1CFE" => data_out<= x"3F";
        when x"1CFF" => data_out<= x"A2";
        when x"1D00" => data_out<= x"B6";
        when x"1D01" => data_out<= x"20";
        when x"1D02" => data_out<= x"F9";
        when x"1D03" => data_out<= x"9A";
        when x"1D04" => data_out<= x"AA";
        when x"1D05" => data_out<= x"F0";
        when x"1D06" => data_out<= x"0E";
        when x"1D07" => data_out<= x"A9";
        when x"1D08" => data_out<= x"0C";
        when x"1D09" => data_out<= x"A2";
        when x"1D0A" => data_out<= x"B6";
        when x"1D0B" => data_out<= x"20";
        when x"1D0C" => data_out<= x"22";
        when x"1D0D" => data_out<= x"81";
        when x"1D0E" => data_out<= x"A9";
        when x"1D0F" => data_out<= x"72";
        when x"1D10" => data_out<= x"A2";
        when x"1D11" => data_out<= x"B3";
        when x"1D12" => data_out<= x"4C";
        when x"1D13" => data_out<= x"F2";
        when x"1D14" => data_out<= x"9D";
        when x"1D15" => data_out<= x"20";
        when x"1D16" => data_out<= x"91";
        when x"1D17" => data_out<= x"B0";
        when x"1D18" => data_out<= x"A9";
        when x"1D19" => data_out<= x"80";
        when x"1D1A" => data_out<= x"A2";
        when x"1D1B" => data_out<= x"BD";
        when x"1D1C" => data_out<= x"20";
        when x"1D1D" => data_out<= x"F9";
        when x"1D1E" => data_out<= x"9A";
        when x"1D1F" => data_out<= x"AA";
        when x"1D20" => data_out<= x"F0";
        when x"1D21" => data_out<= x"0E";
        when x"1D22" => data_out<= x"A9";
        when x"1D23" => data_out<= x"48";
        when x"1D24" => data_out<= x"A2";
        when x"1D25" => data_out<= x"B7";
        when x"1D26" => data_out<= x"20";
        when x"1D27" => data_out<= x"22";
        when x"1D28" => data_out<= x"81";
        when x"1D29" => data_out<= x"A9";
        when x"1D2A" => data_out<= x"C6";
        when x"1D2B" => data_out<= x"A2";
        when x"1D2C" => data_out<= x"B6";
        when x"1D2D" => data_out<= x"4C";
        when x"1D2E" => data_out<= x"F2";
        when x"1D2F" => data_out<= x"9D";
        when x"1D30" => data_out<= x"20";
        when x"1D31" => data_out<= x"91";
        when x"1D32" => data_out<= x"B0";
        when x"1D33" => data_out<= x"A9";
        when x"1D34" => data_out<= x"9A";
        when x"1D35" => data_out<= x"A2";
        when x"1D36" => data_out<= x"BC";
        when x"1D37" => data_out<= x"20";
        when x"1D38" => data_out<= x"F9";
        when x"1D39" => data_out<= x"9A";
        when x"1D3A" => data_out<= x"AA";
        when x"1D3B" => data_out<= x"F0";
        when x"1D3C" => data_out<= x"15";
        when x"1D3D" => data_out<= x"A9";
        when x"1D3E" => data_out<= x"96";
        when x"1D3F" => data_out<= x"A2";
        when x"1D40" => data_out<= x"B9";
        when x"1D41" => data_out<= x"20";
        when x"1D42" => data_out<= x"22";
        when x"1D43" => data_out<= x"81";
        when x"1D44" => data_out<= x"A9";
        when x"1D45" => data_out<= x"3F";
        when x"1D46" => data_out<= x"A2";
        when x"1D47" => data_out<= x"B9";
        when x"1D48" => data_out<= x"20";
        when x"1D49" => data_out<= x"22";
        when x"1D4A" => data_out<= x"81";
        when x"1D4B" => data_out<= x"A9";
        when x"1D4C" => data_out<= x"0B";
        when x"1D4D" => data_out<= x"A2";
        when x"1D4E" => data_out<= x"B5";
        when x"1D4F" => data_out<= x"4C";
        when x"1D50" => data_out<= x"F2";
        when x"1D51" => data_out<= x"9D";
        when x"1D52" => data_out<= x"20";
        when x"1D53" => data_out<= x"91";
        when x"1D54" => data_out<= x"B0";
        when x"1D55" => data_out<= x"A9";
        when x"1D56" => data_out<= x"95";
        when x"1D57" => data_out<= x"A2";
        when x"1D58" => data_out<= x"BC";
        when x"1D59" => data_out<= x"20";
        when x"1D5A" => data_out<= x"F9";
        when x"1D5B" => data_out<= x"9A";
        when x"1D5C" => data_out<= x"AA";
        when x"1D5D" => data_out<= x"F0";
        when x"1D5E" => data_out<= x"1C";
        when x"1D5F" => data_out<= x"A9";
        when x"1D60" => data_out<= x"4B";
        when x"1D61" => data_out<= x"A2";
        when x"1D62" => data_out<= x"BA";
        when x"1D63" => data_out<= x"20";
        when x"1D64" => data_out<= x"22";
        when x"1D65" => data_out<= x"81";
        when x"1D66" => data_out<= x"A9";
        when x"1D67" => data_out<= x"14";
        when x"1D68" => data_out<= x"A2";
        when x"1D69" => data_out<= x"B7";
        when x"1D6A" => data_out<= x"20";
        when x"1D6B" => data_out<= x"22";
        when x"1D6C" => data_out<= x"81";
        when x"1D6D" => data_out<= x"A9";
        when x"1D6E" => data_out<= x"AB";
        when x"1D6F" => data_out<= x"A2";
        when x"1D70" => data_out<= x"B9";
        when x"1D71" => data_out<= x"20";
        when x"1D72" => data_out<= x"22";
        when x"1D73" => data_out<= x"81";
        when x"1D74" => data_out<= x"A9";
        when x"1D75" => data_out<= x"7F";
        when x"1D76" => data_out<= x"A2";
        when x"1D77" => data_out<= x"B2";
        when x"1D78" => data_out<= x"4C";
        when x"1D79" => data_out<= x"F2";
        when x"1D7A" => data_out<= x"9D";
        when x"1D7B" => data_out<= x"20";
        when x"1D7C" => data_out<= x"91";
        when x"1D7D" => data_out<= x"B0";
        when x"1D7E" => data_out<= x"A9";
        when x"1D7F" => data_out<= x"11";
        when x"1D80" => data_out<= x"A2";
        when x"1D81" => data_out<= x"BD";
        when x"1D82" => data_out<= x"20";
        when x"1D83" => data_out<= x"F9";
        when x"1D84" => data_out<= x"9A";
        when x"1D85" => data_out<= x"AA";
        when x"1D86" => data_out<= x"F0";
        when x"1D87" => data_out<= x"0E";
        when x"1D88" => data_out<= x"A9";
        when x"1D89" => data_out<= x"CF";
        when x"1D8A" => data_out<= x"A2";
        when x"1D8B" => data_out<= x"B4";
        when x"1D8C" => data_out<= x"20";
        when x"1D8D" => data_out<= x"22";
        when x"1D8E" => data_out<= x"81";
        when x"1D8F" => data_out<= x"A9";
        when x"1D90" => data_out<= x"10";
        when x"1D91" => data_out<= x"A2";
        when x"1D92" => data_out<= x"BA";
        when x"1D93" => data_out<= x"4C";
        when x"1D94" => data_out<= x"F2";
        when x"1D95" => data_out<= x"9D";
        when x"1D96" => data_out<= x"20";
        when x"1D97" => data_out<= x"91";
        when x"1D98" => data_out<= x"B0";
        when x"1D99" => data_out<= x"A9";
        when x"1D9A" => data_out<= x"39";
        when x"1D9B" => data_out<= x"A2";
        when x"1D9C" => data_out<= x"BD";
        when x"1D9D" => data_out<= x"20";
        when x"1D9E" => data_out<= x"F9";
        when x"1D9F" => data_out<= x"9A";
        when x"1DA0" => data_out<= x"AA";
        when x"1DA1" => data_out<= x"F0";
        when x"1DA2" => data_out<= x"0E";
        when x"1DA3" => data_out<= x"A9";
        when x"1DA4" => data_out<= x"74";
        when x"1DA5" => data_out<= x"A2";
        when x"1DA6" => data_out<= x"B4";
        when x"1DA7" => data_out<= x"20";
        when x"1DA8" => data_out<= x"22";
        when x"1DA9" => data_out<= x"81";
        when x"1DAA" => data_out<= x"A9";
        when x"1DAB" => data_out<= x"38";
        when x"1DAC" => data_out<= x"A2";
        when x"1DAD" => data_out<= x"BA";
        when x"1DAE" => data_out<= x"4C";
        when x"1DAF" => data_out<= x"F2";
        when x"1DB0" => data_out<= x"9D";
        when x"1DB1" => data_out<= x"20";
        when x"1DB2" => data_out<= x"91";
        when x"1DB3" => data_out<= x"B0";
        when x"1DB4" => data_out<= x"A9";
        when x"1DB5" => data_out<= x"0A";
        when x"1DB6" => data_out<= x"A2";
        when x"1DB7" => data_out<= x"BC";
        when x"1DB8" => data_out<= x"20";
        when x"1DB9" => data_out<= x"F9";
        when x"1DBA" => data_out<= x"9A";
        when x"1DBB" => data_out<= x"AA";
        when x"1DBC" => data_out<= x"F0";
        when x"1DBD" => data_out<= x"0E";
        when x"1DBE" => data_out<= x"A9";
        when x"1DBF" => data_out<= x"AC";
        when x"1DC0" => data_out<= x"A2";
        when x"1DC1" => data_out<= x"B6";
        when x"1DC2" => data_out<= x"20";
        when x"1DC3" => data_out<= x"22";
        when x"1DC4" => data_out<= x"81";
        when x"1DC5" => data_out<= x"A9";
        when x"1DC6" => data_out<= x"D5";
        when x"1DC7" => data_out<= x"A2";
        when x"1DC8" => data_out<= x"B5";
        when x"1DC9" => data_out<= x"4C";
        when x"1DCA" => data_out<= x"F2";
        when x"1DCB" => data_out<= x"9D";
        when x"1DCC" => data_out<= x"20";
        when x"1DCD" => data_out<= x"91";
        when x"1DCE" => data_out<= x"B0";
        when x"1DCF" => data_out<= x"A9";
        when x"1DD0" => data_out<= x"61";
        when x"1DD1" => data_out<= x"A2";
        when x"1DD2" => data_out<= x"BC";
        when x"1DD3" => data_out<= x"20";
        when x"1DD4" => data_out<= x"F9";
        when x"1DD5" => data_out<= x"9A";
        when x"1DD6" => data_out<= x"AA";
        when x"1DD7" => data_out<= x"F0";
        when x"1DD8" => data_out<= x"15";
        when x"1DD9" => data_out<= x"A9";
        when x"1DDA" => data_out<= x"35";
        when x"1DDB" => data_out<= x"A2";
        when x"1DDC" => data_out<= x"B4";
        when x"1DDD" => data_out<= x"20";
        when x"1DDE" => data_out<= x"22";
        when x"1DDF" => data_out<= x"81";
        when x"1DE0" => data_out<= x"A9";
        when x"1DE1" => data_out<= x"AB";
        when x"1DE2" => data_out<= x"A2";
        when x"1DE3" => data_out<= x"B9";
        when x"1DE4" => data_out<= x"20";
        when x"1DE5" => data_out<= x"22";
        when x"1DE6" => data_out<= x"81";
        when x"1DE7" => data_out<= x"A9";
        when x"1DE8" => data_out<= x"6E";
        when x"1DE9" => data_out<= x"A2";
        when x"1DEA" => data_out<= x"B8";
        when x"1DEB" => data_out<= x"4C";
        when x"1DEC" => data_out<= x"F2";
        when x"1DED" => data_out<= x"9D";
        when x"1DEE" => data_out<= x"A9";
        when x"1DEF" => data_out<= x"E1";
        when x"1DF0" => data_out<= x"A2";
        when x"1DF1" => data_out<= x"B1";
        when x"1DF2" => data_out<= x"20";
        when x"1DF3" => data_out<= x"22";
        when x"1DF4" => data_out<= x"81";
        when x"1DF5" => data_out<= x"4C";
        when x"1DF6" => data_out<= x"14";
        when x"1DF7" => data_out<= x"AF";
        when x"1DF8" => data_out<= x"20";
        when x"1DF9" => data_out<= x"65";
        when x"1DFA" => data_out<= x"B0";
        when x"1DFB" => data_out<= x"A9";
        when x"1DFC" => data_out<= x"00";
        when x"1DFD" => data_out<= x"20";
        when x"1DFE" => data_out<= x"65";
        when x"1DFF" => data_out<= x"B0";
        when x"1E00" => data_out<= x"20";
        when x"1E01" => data_out<= x"6A";
        when x"1E02" => data_out<= x"AE";
        when x"1E03" => data_out<= x"4C";
        when x"1E04" => data_out<= x"13";
        when x"1E05" => data_out<= x"9E";
        when x"1E06" => data_out<= x"A0";
        when x"1E07" => data_out<= x"06";
        when x"1E08" => data_out<= x"20";
        when x"1E09" => data_out<= x"4F";
        when x"1E0A" => data_out<= x"AF";
        when x"1E0B" => data_out<= x"20";
        when x"1E0C" => data_out<= x"E2";
        when x"1E0D" => data_out<= x"AE";
        when x"1E0E" => data_out<= x"A0";
        when x"1E0F" => data_out<= x"05";
        when x"1E10" => data_out<= x"20";
        when x"1E11" => data_out<= x"C5";
        when x"1E12" => data_out<= x"B0";
        when x"1E13" => data_out<= x"A0";
        when x"1E14" => data_out<= x"06";
        when x"1E15" => data_out<= x"20";
        when x"1E16" => data_out<= x"4F";
        when x"1E17" => data_out<= x"AF";
        when x"1E18" => data_out<= x"85";
        when x"1E19" => data_out<= x"14";
        when x"1E1A" => data_out<= x"86";
        when x"1E1B" => data_out<= x"15";
        when x"1E1C" => data_out<= x"A0";
        when x"1E1D" => data_out<= x"00";
        when x"1E1E" => data_out<= x"B1";
        when x"1E1F" => data_out<= x"14";
        when x"1E20" => data_out<= x"C9";
        when x"1E21" => data_out<= x"20";
        when x"1E22" => data_out<= x"F0";
        when x"1E23" => data_out<= x"E2";
        when x"1E24" => data_out<= x"4C";
        when x"1E25" => data_out<= x"6A";
        when x"1E26" => data_out<= x"9E";
        when x"1E27" => data_out<= x"A0";
        when x"1E28" => data_out<= x"06";
        when x"1E29" => data_out<= x"20";
        when x"1E2A" => data_out<= x"4F";
        when x"1E2B" => data_out<= x"AF";
        when x"1E2C" => data_out<= x"85";
        when x"1E2D" => data_out<= x"10";
        when x"1E2E" => data_out<= x"86";
        when x"1E2F" => data_out<= x"11";
        when x"1E30" => data_out<= x"20";
        when x"1E31" => data_out<= x"E2";
        when x"1E32" => data_out<= x"AE";
        when x"1E33" => data_out<= x"A0";
        when x"1E34" => data_out<= x"05";
        when x"1E35" => data_out<= x"20";
        when x"1E36" => data_out<= x"C5";
        when x"1E37" => data_out<= x"B0";
        when x"1E38" => data_out<= x"A0";
        when x"1E39" => data_out<= x"00";
        when x"1E3A" => data_out<= x"B1";
        when x"1E3B" => data_out<= x"10";
        when x"1E3C" => data_out<= x"91";
        when x"1E3D" => data_out<= x"0C";
        when x"1E3E" => data_out<= x"C9";
        when x"1E3F" => data_out<= x"61";
        when x"1E40" => data_out<= x"90";
        when x"1E41" => data_out<= x"0B";
        when x"1E42" => data_out<= x"B1";
        when x"1E43" => data_out<= x"0C";
        when x"1E44" => data_out<= x"C9";
        when x"1E45" => data_out<= x"7B";
        when x"1E46" => data_out<= x"B0";
        when x"1E47" => data_out<= x"05";
        when x"1E48" => data_out<= x"38";
        when x"1E49" => data_out<= x"E9";
        when x"1E4A" => data_out<= x"20";
        when x"1E4B" => data_out<= x"91";
        when x"1E4C" => data_out<= x"0C";
        when x"1E4D" => data_out<= x"A0";
        when x"1E4E" => data_out<= x"06";
        when x"1E4F" => data_out<= x"20";
        when x"1E50" => data_out<= x"93";
        when x"1E51" => data_out<= x"B0";
        when x"1E52" => data_out<= x"A0";
        when x"1E53" => data_out<= x"03";
        when x"1E54" => data_out<= x"B1";
        when x"1E55" => data_out<= x"0C";
        when x"1E56" => data_out<= x"48";
        when x"1E57" => data_out<= x"18";
        when x"1E58" => data_out<= x"69";
        when x"1E59" => data_out<= x"01";
        when x"1E5A" => data_out<= x"91";
        when x"1E5B" => data_out<= x"0C";
        when x"1E5C" => data_out<= x"68";
        when x"1E5D" => data_out<= x"20";
        when x"1E5E" => data_out<= x"E6";
        when x"1E5F" => data_out<= x"AD";
        when x"1E60" => data_out<= x"85";
        when x"1E61" => data_out<= x"14";
        when x"1E62" => data_out<= x"86";
        when x"1E63" => data_out<= x"15";
        when x"1E64" => data_out<= x"A0";
        when x"1E65" => data_out<= x"00";
        when x"1E66" => data_out<= x"B1";
        when x"1E67" => data_out<= x"0C";
        when x"1E68" => data_out<= x"91";
        when x"1E69" => data_out<= x"14";
        when x"1E6A" => data_out<= x"A0";
        when x"1E6B" => data_out<= x"06";
        when x"1E6C" => data_out<= x"20";
        when x"1E6D" => data_out<= x"4F";
        when x"1E6E" => data_out<= x"AF";
        when x"1E6F" => data_out<= x"85";
        when x"1E70" => data_out<= x"14";
        when x"1E71" => data_out<= x"86";
        when x"1E72" => data_out<= x"15";
        when x"1E73" => data_out<= x"A0";
        when x"1E74" => data_out<= x"00";
        when x"1E75" => data_out<= x"B1";
        when x"1E76" => data_out<= x"14";
        when x"1E77" => data_out<= x"F0";
        when x"1E78" => data_out<= x"23";
        when x"1E79" => data_out<= x"A0";
        when x"1E7A" => data_out<= x"06";
        when x"1E7B" => data_out<= x"20";
        when x"1E7C" => data_out<= x"4F";
        when x"1E7D" => data_out<= x"AF";
        when x"1E7E" => data_out<= x"85";
        when x"1E7F" => data_out<= x"14";
        when x"1E80" => data_out<= x"86";
        when x"1E81" => data_out<= x"15";
        when x"1E82" => data_out<= x"A0";
        when x"1E83" => data_out<= x"00";
        when x"1E84" => data_out<= x"B1";
        when x"1E85" => data_out<= x"14";
        when x"1E86" => data_out<= x"C9";
        when x"1E87" => data_out<= x"20";
        when x"1E88" => data_out<= x"F0";
        when x"1E89" => data_out<= x"12";
        when x"1E8A" => data_out<= x"C8";
        when x"1E8B" => data_out<= x"B1";
        when x"1E8C" => data_out<= x"0C";
        when x"1E8D" => data_out<= x"20";
        when x"1E8E" => data_out<= x"79";
        when x"1E8F" => data_out<= x"B0";
        when x"1E90" => data_out<= x"A0";
        when x"1E91" => data_out<= x"04";
        when x"1E92" => data_out<= x"B1";
        when x"1E93" => data_out<= x"0C";
        when x"1E94" => data_out<= x"20";
        when x"1E95" => data_out<= x"5A";
        when x"1E96" => data_out<= x"AE";
        when x"1E97" => data_out<= x"20";
        when x"1E98" => data_out<= x"B6";
        when x"1E99" => data_out<= x"AE";
        when x"1E9A" => data_out<= x"90";
        when x"1E9B" => data_out<= x"8B";
        when x"1E9C" => data_out<= x"A0";
        when x"1E9D" => data_out<= x"01";
        when x"1E9E" => data_out<= x"B1";
        when x"1E9F" => data_out<= x"0C";
        when x"1EA0" => data_out<= x"18";
        when x"1EA1" => data_out<= x"A0";
        when x"1EA2" => data_out<= x"03";
        when x"1EA3" => data_out<= x"71";
        when x"1EA4" => data_out<= x"0C";
        when x"1EA5" => data_out<= x"85";
        when x"1EA6" => data_out<= x"14";
        when x"1EA7" => data_out<= x"A9";
        when x"1EA8" => data_out<= x"00";
        when x"1EA9" => data_out<= x"C8";
        when x"1EAA" => data_out<= x"71";
        when x"1EAB" => data_out<= x"0C";
        when x"1EAC" => data_out<= x"85";
        when x"1EAD" => data_out<= x"15";
        when x"1EAE" => data_out<= x"A9";
        when x"1EAF" => data_out<= x"00";
        when x"1EB0" => data_out<= x"A8";
        when x"1EB1" => data_out<= x"91";
        when x"1EB2" => data_out<= x"14";
        when x"1EB3" => data_out<= x"A0";
        when x"1EB4" => data_out<= x"06";
        when x"1EB5" => data_out<= x"20";
        when x"1EB6" => data_out<= x"4F";
        when x"1EB7" => data_out<= x"AF";
        when x"1EB8" => data_out<= x"4C";
        when x"1EB9" => data_out<= x"36";
        when x"1EBA" => data_out<= x"AF";
        when x"1EBB" => data_out<= x"20";
        when x"1EBC" => data_out<= x"6A";
        when x"1EBD" => data_out<= x"AE";
        when x"1EBE" => data_out<= x"A9";
        when x"1EBF" => data_out<= x"00";
        when x"1EC0" => data_out<= x"8D";
        when x"1EC1" => data_out<= x"46";
        when x"1EC2" => data_out<= x"02";
        when x"1EC3" => data_out<= x"20";
        when x"1EC4" => data_out<= x"FD";
        when x"1EC5" => data_out<= x"80";
        when x"1EC6" => data_out<= x"A0";
        when x"1EC7" => data_out<= x"00";
        when x"1EC8" => data_out<= x"91";
        when x"1EC9" => data_out<= x"0C";
        when x"1ECA" => data_out<= x"C9";
        when x"1ECB" => data_out<= x"0D";
        when x"1ECC" => data_out<= x"F0";
        when x"1ECD" => data_out<= x"06";
        when x"1ECE" => data_out<= x"B1";
        when x"1ECF" => data_out<= x"0C";
        when x"1ED0" => data_out<= x"C9";
        when x"1ED1" => data_out<= x"0A";
        when x"1ED2" => data_out<= x"D0";
        when x"1ED3" => data_out<= x"0E";
        when x"1ED4" => data_out<= x"AC";
        when x"1ED5" => data_out<= x"46";
        when x"1ED6" => data_out<= x"02";
        when x"1ED7" => data_out<= x"A9";
        when x"1ED8" => data_out<= x"00";
        when x"1ED9" => data_out<= x"99";
        when x"1EDA" => data_out<= x"06";
        when x"1EDB" => data_out<= x"02";
        when x"1EDC" => data_out<= x"20";
        when x"1EDD" => data_out<= x"45";
        when x"1EDE" => data_out<= x"8C";
        when x"1EDF" => data_out<= x"4C";
        when x"1EE0" => data_out<= x"05";
        when x"1EE1" => data_out<= x"AF";
        when x"1EE2" => data_out<= x"B1";
        when x"1EE3" => data_out<= x"0C";
        when x"1EE4" => data_out<= x"C9";
        when x"1EE5" => data_out<= x"08";
        when x"1EE6" => data_out<= x"F0";
        when x"1EE7" => data_out<= x"04";
        when x"1EE8" => data_out<= x"C9";
        when x"1EE9" => data_out<= x"7F";
        when x"1EEA" => data_out<= x"D0";
        when x"1EEB" => data_out<= x"1A";
        when x"1EEC" => data_out<= x"AD";
        when x"1EED" => data_out<= x"46";
        when x"1EEE" => data_out<= x"02";
        when x"1EEF" => data_out<= x"F0";
        when x"1EF0" => data_out<= x"D2";
        when x"1EF1" => data_out<= x"CE";
        when x"1EF2" => data_out<= x"46";
        when x"1EF3" => data_out<= x"02";
        when x"1EF4" => data_out<= x"A9";
        when x"1EF5" => data_out<= x"08";
        when x"1EF6" => data_out<= x"20";
        when x"1EF7" => data_out<= x"F0";
        when x"1EF8" => data_out<= x"80";
        when x"1EF9" => data_out<= x"A9";
        when x"1EFA" => data_out<= x"20";
        when x"1EFB" => data_out<= x"20";
        when x"1EFC" => data_out<= x"F0";
        when x"1EFD" => data_out<= x"80";
        when x"1EFE" => data_out<= x"A9";
        when x"1EFF" => data_out<= x"08";
        when x"1F00" => data_out<= x"20";
        when x"1F01" => data_out<= x"F0";
        when x"1F02" => data_out<= x"80";
        when x"1F03" => data_out<= x"4C";
        when x"1F04" => data_out<= x"C3";
        when x"1F05" => data_out<= x"9E";
        when x"1F06" => data_out<= x"B1";
        when x"1F07" => data_out<= x"0C";
        when x"1F08" => data_out<= x"C9";
        when x"1F09" => data_out<= x"1B";
        when x"1F0A" => data_out<= x"D0";
        when x"1F0B" => data_out<= x"14";
        when x"1F0C" => data_out<= x"98";
        when x"1F0D" => data_out<= x"8D";
        when x"1F0E" => data_out<= x"46";
        when x"1F0F" => data_out<= x"02";
        when x"1F10" => data_out<= x"8D";
        when x"1F11" => data_out<= x"06";
        when x"1F12" => data_out<= x"02";
        when x"1F13" => data_out<= x"A9";
        when x"1F14" => data_out<= x"3B";
        when x"1F15" => data_out<= x"A2";
        when x"1F16" => data_out<= x"BC";
        when x"1F17" => data_out<= x"20";
        when x"1F18" => data_out<= x"22";
        when x"1F19" => data_out<= x"81";
        when x"1F1A" => data_out<= x"20";
        when x"1F1B" => data_out<= x"45";
        when x"1F1C" => data_out<= x"8C";
        when x"1F1D" => data_out<= x"4C";
        when x"1F1E" => data_out<= x"05";
        when x"1F1F" => data_out<= x"AF";
        when x"1F20" => data_out<= x"AD";
        when x"1F21" => data_out<= x"46";
        when x"1F22" => data_out<= x"02";
        when x"1F23" => data_out<= x"C9";
        when x"1F24" => data_out<= x"3F";
        when x"1F25" => data_out<= x"B0";
        when x"1F26" => data_out<= x"9C";
        when x"1F27" => data_out<= x"B1";
        when x"1F28" => data_out<= x"0C";
        when x"1F29" => data_out<= x"C9";
        when x"1F2A" => data_out<= x"20";
        when x"1F2B" => data_out<= x"90";
        when x"1F2C" => data_out<= x"96";
        when x"1F2D" => data_out<= x"C9";
        when x"1F2E" => data_out<= x"7F";
        when x"1F2F" => data_out<= x"B0";
        when x"1F30" => data_out<= x"92";
        when x"1F31" => data_out<= x"AD";
        when x"1F32" => data_out<= x"46";
        when x"1F33" => data_out<= x"02";
        when x"1F34" => data_out<= x"EE";
        when x"1F35" => data_out<= x"46";
        when x"1F36" => data_out<= x"02";
        when x"1F37" => data_out<= x"18";
        when x"1F38" => data_out<= x"69";
        when x"1F39" => data_out<= x"06";
        when x"1F3A" => data_out<= x"85";
        when x"1F3B" => data_out<= x"14";
        when x"1F3C" => data_out<= x"98";
        when x"1F3D" => data_out<= x"69";
        when x"1F3E" => data_out<= x"02";
        when x"1F3F" => data_out<= x"85";
        when x"1F40" => data_out<= x"15";
        when x"1F41" => data_out<= x"B1";
        when x"1F42" => data_out<= x"0C";
        when x"1F43" => data_out<= x"91";
        when x"1F44" => data_out<= x"14";
        when x"1F45" => data_out<= x"B1";
        when x"1F46" => data_out<= x"0C";
        when x"1F47" => data_out<= x"20";
        when x"1F48" => data_out<= x"F0";
        when x"1F49" => data_out<= x"80";
        when x"1F4A" => data_out<= x"4C";
        when x"1F4B" => data_out<= x"C3";
        when x"1F4C" => data_out<= x"9E";
        when x"1F4D" => data_out<= x"A9";
        when x"1F4E" => data_out<= x"00";
        when x"1F4F" => data_out<= x"8D";
        when x"1F50" => data_out<= x"44";
        when x"1F51" => data_out<= x"C0";
        when x"1F52" => data_out<= x"8D";
        when x"1F53" => data_out<= x"45";
        when x"1F54" => data_out<= x"C0";
        when x"1F55" => data_out<= x"60";
        when x"1F56" => data_out<= x"8D";
        when x"1F57" => data_out<= x"44";
        when x"1F58" => data_out<= x"C0";
        when x"1F59" => data_out<= x"A9";
        when x"1F5A" => data_out<= x"01";
        when x"1F5B" => data_out<= x"8D";
        when x"1F5C" => data_out<= x"45";
        when x"1F5D" => data_out<= x"C0";
        when x"1F5E" => data_out<= x"60";
        when x"1F5F" => data_out<= x"A9";
        when x"1F60" => data_out<= x"00";
        when x"1F61" => data_out<= x"8D";
        when x"1F62" => data_out<= x"45";
        when x"1F63" => data_out<= x"C0";
        when x"1F64" => data_out<= x"60";
        when x"1F65" => data_out<= x"48";
        when x"1F66" => data_out<= x"AD";
        when x"1F67" => data_out<= x"42";
        when x"1F68" => data_out<= x"C0";
        when x"1F69" => data_out<= x"29";
        when x"1F6A" => data_out<= x"20";
        when x"1F6B" => data_out<= x"F0";
        when x"1F6C" => data_out<= x"F9";
        when x"1F6D" => data_out<= x"68";
        when x"1F6E" => data_out<= x"8D";
        when x"1F6F" => data_out<= x"41";
        when x"1F70" => data_out<= x"C0";
        when x"1F71" => data_out<= x"AD";
        when x"1F72" => data_out<= x"42";
        when x"1F73" => data_out<= x"C0";
        when x"1F74" => data_out<= x"29";
        when x"1F75" => data_out<= x"40";
        when x"1F76" => data_out<= x"F0";
        when x"1F77" => data_out<= x"F9";
        when x"1F78" => data_out<= x"AD";
        when x"1F79" => data_out<= x"40";
        when x"1F7A" => data_out<= x"C0";
        when x"1F7B" => data_out<= x"A2";
        when x"1F7C" => data_out<= x"00";
        when x"1F7D" => data_out<= x"60";
        when x"1F7E" => data_out<= x"48";
        when x"1F7F" => data_out<= x"AD";
        when x"1F80" => data_out<= x"42";
        when x"1F81" => data_out<= x"C0";
        when x"1F82" => data_out<= x"29";
        when x"1F83" => data_out<= x"20";
        when x"1F84" => data_out<= x"F0";
        when x"1F85" => data_out<= x"F9";
        when x"1F86" => data_out<= x"68";
        when x"1F87" => data_out<= x"8D";
        when x"1F88" => data_out<= x"41";
        when x"1F89" => data_out<= x"C0";
        when x"1F8A" => data_out<= x"AD";
        when x"1F8B" => data_out<= x"42";
        when x"1F8C" => data_out<= x"C0";
        when x"1F8D" => data_out<= x"29";
        when x"1F8E" => data_out<= x"40";
        when x"1F8F" => data_out<= x"F0";
        when x"1F90" => data_out<= x"F9";
        when x"1F91" => data_out<= x"AD";
        when x"1F92" => data_out<= x"40";
        when x"1F93" => data_out<= x"C0";
        when x"1F94" => data_out<= x"60";
        when x"1F95" => data_out<= x"AD";
        when x"1F96" => data_out<= x"42";
        when x"1F97" => data_out<= x"C0";
        when x"1F98" => data_out<= x"29";
        when x"1F99" => data_out<= x"20";
        when x"1F9A" => data_out<= x"F0";
        when x"1F9B" => data_out<= x"F9";
        when x"1F9C" => data_out<= x"A9";
        when x"1F9D" => data_out<= x"FF";
        when x"1F9E" => data_out<= x"8D";
        when x"1F9F" => data_out<= x"41";
        when x"1FA0" => data_out<= x"C0";
        when x"1FA1" => data_out<= x"AD";
        when x"1FA2" => data_out<= x"42";
        when x"1FA3" => data_out<= x"C0";
        when x"1FA4" => data_out<= x"29";
        when x"1FA5" => data_out<= x"40";
        when x"1FA6" => data_out<= x"F0";
        when x"1FA7" => data_out<= x"F9";
        when x"1FA8" => data_out<= x"AD";
        when x"1FA9" => data_out<= x"40";
        when x"1FAA" => data_out<= x"C0";
        when x"1FAB" => data_out<= x"A2";
        when x"1FAC" => data_out<= x"00";
        when x"1FAD" => data_out<= x"60";
        when x"1FAE" => data_out<= x"AD";
        when x"1FAF" => data_out<= x"42";
        when x"1FB0" => data_out<= x"C0";
        when x"1FB1" => data_out<= x"29";
        when x"1FB2" => data_out<= x"20";
        when x"1FB3" => data_out<= x"F0";
        when x"1FB4" => data_out<= x"05";
        when x"1FB5" => data_out<= x"A9";
        when x"1FB6" => data_out<= x"00";
        when x"1FB7" => data_out<= x"A2";
        when x"1FB8" => data_out<= x"00";
        when x"1FB9" => data_out<= x"60";
        when x"1FBA" => data_out<= x"A9";
        when x"1FBB" => data_out<= x"01";
        when x"1FBC" => data_out<= x"A2";
        when x"1FBD" => data_out<= x"00";
        when x"1FBE" => data_out<= x"60";
        when x"1FBF" => data_out<= x"20";
        when x"1FC0" => data_out<= x"8D";
        when x"1FC1" => data_out<= x"AE";
        when x"1FC2" => data_out<= x"A9";
        when x"1FC3" => data_out<= x"00";
        when x"1FC4" => data_out<= x"8D";
        when x"1FC5" => data_out<= x"05";
        when x"1FC6" => data_out<= x"02";
        when x"1FC7" => data_out<= x"8D";
        when x"1FC8" => data_out<= x"04";
        when x"1FC9" => data_out<= x"02";
        when x"1FCA" => data_out<= x"20";
        when x"1FCB" => data_out<= x"4D";
        when x"1FCC" => data_out<= x"9F";
        when x"1FCD" => data_out<= x"20";
        when x"1FCE" => data_out<= x"7C";
        when x"1FCF" => data_out<= x"A2";
        when x"1FD0" => data_out<= x"A9";
        when x"1FD1" => data_out<= x"00";
        when x"1FD2" => data_out<= x"A0";
        when x"1FD3" => data_out<= x"02";
        when x"1FD4" => data_out<= x"91";
        when x"1FD5" => data_out<= x"0C";
        when x"1FD6" => data_out<= x"C9";
        when x"1FD7" => data_out<= x"0A";
        when x"1FD8" => data_out<= x"B0";
        when x"1FD9" => data_out<= x"0F";
        when x"1FDA" => data_out<= x"A9";
        when x"1FDB" => data_out<= x"FF";
        when x"1FDC" => data_out<= x"20";
        when x"1FDD" => data_out<= x"65";
        when x"1FDE" => data_out<= x"9F";
        when x"1FDF" => data_out<= x"A0";
        when x"1FE0" => data_out<= x"02";
        when x"1FE1" => data_out<= x"B1";
        when x"1FE2" => data_out<= x"0C";
        when x"1FE3" => data_out<= x"18";
        when x"1FE4" => data_out<= x"69";
        when x"1FE5" => data_out<= x"01";
        when x"1FE6" => data_out<= x"4C";
        when x"1FE7" => data_out<= x"D4";
        when x"1FE8" => data_out<= x"9F";
        when x"1FE9" => data_out<= x"20";
        when x"1FEA" => data_out<= x"77";
        when x"1FEB" => data_out<= x"A2";
        when x"1FEC" => data_out<= x"A9";
        when x"1FED" => data_out<= x"40";
        when x"1FEE" => data_out<= x"20";
        when x"1FEF" => data_out<= x"65";
        when x"1FF0" => data_out<= x"B0";
        when x"1FF1" => data_out<= x"20";
        when x"1FF2" => data_out<= x"75";
        when x"1FF3" => data_out<= x"AF";
        when x"1FF4" => data_out<= x"A9";
        when x"1FF5" => data_out<= x"95";
        when x"1FF6" => data_out<= x"20";
        when x"1FF7" => data_out<= x"7F";
        when x"1FF8" => data_out<= x"A2";
        when x"1FF9" => data_out<= x"A0";
        when x"1FFA" => data_out<= x"03";
        when x"1FFB" => data_out<= x"91";
        when x"1FFC" => data_out<= x"0C";
        when x"1FFD" => data_out<= x"20";
        when x"1FFE" => data_out<= x"7C";
        when x"1FFF" => data_out<= x"A2";
        when x"2000" => data_out<= x"A9";
        when x"2001" => data_out<= x"FF";
        when x"2002" => data_out<= x"20";
        when x"2003" => data_out<= x"65";
        when x"2004" => data_out<= x"9F";
        when x"2005" => data_out<= x"A0";
        when x"2006" => data_out<= x"03";
        when x"2007" => data_out<= x"B1";
        when x"2008" => data_out<= x"0C";
        when x"2009" => data_out<= x"C9";
        when x"200A" => data_out<= x"01";
        when x"200B" => data_out<= x"F0";
        when x"200C" => data_out<= x"06";
        when x"200D" => data_out<= x"A2";
        when x"200E" => data_out<= x"00";
        when x"200F" => data_out<= x"98";
        when x"2010" => data_out<= x"4C";
        when x"2011" => data_out<= x"27";
        when x"2012" => data_out<= x"AF";
        when x"2013" => data_out<= x"20";
        when x"2014" => data_out<= x"77";
        when x"2015" => data_out<= x"A2";
        when x"2016" => data_out<= x"A9";
        when x"2017" => data_out<= x"48";
        when x"2018" => data_out<= x"20";
        when x"2019" => data_out<= x"65";
        when x"201A" => data_out<= x"B0";
        when x"201B" => data_out<= x"A2";
        when x"201C" => data_out<= x"01";
        when x"201D" => data_out<= x"A9";
        when x"201E" => data_out<= x"AA";
        when x"201F" => data_out<= x"20";
        when x"2020" => data_out<= x"78";
        when x"2021" => data_out<= x"AF";
        when x"2022" => data_out<= x"A9";
        when x"2023" => data_out<= x"87";
        when x"2024" => data_out<= x"20";
        when x"2025" => data_out<= x"7F";
        when x"2026" => data_out<= x"A2";
        when x"2027" => data_out<= x"A0";
        when x"2028" => data_out<= x"03";
        when x"2029" => data_out<= x"91";
        when x"202A" => data_out<= x"0C";
        when x"202B" => data_out<= x"C9";
        when x"202C" => data_out<= x"01";
        when x"202D" => data_out<= x"D0";
        when x"202E" => data_out<= x"19";
        when x"202F" => data_out<= x"A9";
        when x"2030" => data_out<= x"FF";
        when x"2031" => data_out<= x"20";
        when x"2032" => data_out<= x"65";
        when x"2033" => data_out<= x"9F";
        when x"2034" => data_out<= x"A9";
        when x"2035" => data_out<= x"FF";
        when x"2036" => data_out<= x"20";
        when x"2037" => data_out<= x"65";
        when x"2038" => data_out<= x"9F";
        when x"2039" => data_out<= x"A9";
        when x"203A" => data_out<= x"FF";
        when x"203B" => data_out<= x"20";
        when x"203C" => data_out<= x"65";
        when x"203D" => data_out<= x"9F";
        when x"203E" => data_out<= x"A9";
        when x"203F" => data_out<= x"FF";
        when x"2040" => data_out<= x"20";
        when x"2041" => data_out<= x"65";
        when x"2042" => data_out<= x"9F";
        when x"2043" => data_out<= x"A9";
        when x"2044" => data_out<= x"02";
        when x"2045" => data_out<= x"4C";
        when x"2046" => data_out<= x"4A";
        when x"2047" => data_out<= x"A0";
        when x"2048" => data_out<= x"A9";
        when x"2049" => data_out<= x"01";
        when x"204A" => data_out<= x"8D";
        when x"204B" => data_out<= x"04";
        when x"204C" => data_out<= x"02";
        when x"204D" => data_out<= x"20";
        when x"204E" => data_out<= x"7C";
        when x"204F" => data_out<= x"A2";
        when x"2050" => data_out<= x"A9";
        when x"2051" => data_out<= x"FF";
        when x"2052" => data_out<= x"20";
        when x"2053" => data_out<= x"65";
        when x"2054" => data_out<= x"9F";
        when x"2055" => data_out<= x"A2";
        when x"2056" => data_out<= x"00";
        when x"2057" => data_out<= x"8A";
        when x"2058" => data_out<= x"20";
        when x"2059" => data_out<= x"C3";
        when x"205A" => data_out<= x"B0";
        when x"205B" => data_out<= x"A0";
        when x"205C" => data_out<= x"01";
        when x"205D" => data_out<= x"B1";
        when x"205E" => data_out<= x"0C";
        when x"205F" => data_out<= x"C9";
        when x"2060" => data_out<= x"03";
        when x"2061" => data_out<= x"D0";
        when x"2062" => data_out<= x"05";
        when x"2063" => data_out<= x"88";
        when x"2064" => data_out<= x"B1";
        when x"2065" => data_out<= x"0C";
        when x"2066" => data_out<= x"C9";
        when x"2067" => data_out<= x"E8";
        when x"2068" => data_out<= x"B0";
        when x"2069" => data_out<= x"3D";
        when x"206A" => data_out<= x"20";
        when x"206B" => data_out<= x"77";
        when x"206C" => data_out<= x"A2";
        when x"206D" => data_out<= x"A9";
        when x"206E" => data_out<= x"69";
        when x"206F" => data_out<= x"20";
        when x"2070" => data_out<= x"65";
        when x"2071" => data_out<= x"B0";
        when x"2072" => data_out<= x"A2";
        when x"2073" => data_out<= x"00";
        when x"2074" => data_out<= x"AD";
        when x"2075" => data_out<= x"04";
        when x"2076" => data_out<= x"02";
        when x"2077" => data_out<= x"C9";
        when x"2078" => data_out<= x"02";
        when x"2079" => data_out<= x"D0";
        when x"207A" => data_out<= x"0A";
        when x"207B" => data_out<= x"86";
        when x"207C" => data_out<= x"0E";
        when x"207D" => data_out<= x"A9";
        when x"207E" => data_out<= x"40";
        when x"207F" => data_out<= x"85";
        when x"2080" => data_out<= x"0F";
        when x"2081" => data_out<= x"8A";
        when x"2082" => data_out<= x"4C";
        when x"2083" => data_out<= x"89";
        when x"2084" => data_out<= x"A0";
        when x"2085" => data_out<= x"8A";
        when x"2086" => data_out<= x"20";
        when x"2087" => data_out<= x"46";
        when x"2088" => data_out<= x"AE";
        when x"2089" => data_out<= x"20";
        when x"208A" => data_out<= x"EF";
        when x"208B" => data_out<= x"A2";
        when x"208C" => data_out<= x"A0";
        when x"208D" => data_out<= x"03";
        when x"208E" => data_out<= x"91";
        when x"208F" => data_out<= x"0C";
        when x"2090" => data_out<= x"20";
        when x"2091" => data_out<= x"7C";
        when x"2092" => data_out<= x"A2";
        when x"2093" => data_out<= x"A9";
        when x"2094" => data_out<= x"FF";
        when x"2095" => data_out<= x"20";
        when x"2096" => data_out<= x"65";
        when x"2097" => data_out<= x"9F";
        when x"2098" => data_out<= x"A0";
        when x"2099" => data_out<= x"03";
        when x"209A" => data_out<= x"B1";
        when x"209B" => data_out<= x"0C";
        when x"209C" => data_out<= x"F0";
        when x"209D" => data_out<= x"0B";
        when x"209E" => data_out<= x"20";
        when x"209F" => data_out<= x"4D";
        when x"20A0" => data_out<= x"AF";
        when x"20A1" => data_out<= x"20";
        when x"20A2" => data_out<= x"E2";
        when x"20A3" => data_out<= x"AE";
        when x"20A4" => data_out<= x"4C";
        when x"20A5" => data_out<= x"58";
        when x"20A6" => data_out<= x"A0";
        when x"20A7" => data_out<= x"A0";
        when x"20A8" => data_out<= x"03";
        when x"20A9" => data_out<= x"B1";
        when x"20AA" => data_out<= x"0C";
        when x"20AB" => data_out<= x"F0";
        when x"20AC" => data_out<= x"07";
        when x"20AD" => data_out<= x"A2";
        when x"20AE" => data_out<= x"00";
        when x"20AF" => data_out<= x"A9";
        when x"20B0" => data_out<= x"01";
        when x"20B1" => data_out<= x"4C";
        when x"20B2" => data_out<= x"27";
        when x"20B3" => data_out<= x"AF";
        when x"20B4" => data_out<= x"AD";
        when x"20B5" => data_out<= x"04";
        when x"20B6" => data_out<= x"02";
        when x"20B7" => data_out<= x"C9";
        when x"20B8" => data_out<= x"02";
        when x"20B9" => data_out<= x"D0";
        when x"20BA" => data_out<= x"47";
        when x"20BB" => data_out<= x"20";
        when x"20BC" => data_out<= x"77";
        when x"20BD" => data_out<= x"A2";
        when x"20BE" => data_out<= x"A9";
        when x"20BF" => data_out<= x"7A";
        when x"20C0" => data_out<= x"20";
        when x"20C1" => data_out<= x"65";
        when x"20C2" => data_out<= x"B0";
        when x"20C3" => data_out<= x"20";
        when x"20C4" => data_out<= x"75";
        when x"20C5" => data_out<= x"AF";
        when x"20C6" => data_out<= x"A9";
        when x"20C7" => data_out<= x"FF";
        when x"20C8" => data_out<= x"20";
        when x"20C9" => data_out<= x"7F";
        when x"20CA" => data_out<= x"A2";
        when x"20CB" => data_out<= x"A0";
        when x"20CC" => data_out<= x"03";
        when x"20CD" => data_out<= x"91";
        when x"20CE" => data_out<= x"0C";
        when x"20CF" => data_out<= x"B1";
        when x"20D0" => data_out<= x"0C";
        when x"20D1" => data_out<= x"D0";
        when x"20D2" => data_out<= x"27";
        when x"20D3" => data_out<= x"A9";
        when x"20D4" => data_out<= x"FF";
        when x"20D5" => data_out<= x"20";
        when x"20D6" => data_out<= x"65";
        when x"20D7" => data_out<= x"9F";
        when x"20D8" => data_out<= x"20";
        when x"20D9" => data_out<= x"65";
        when x"20DA" => data_out<= x"B0";
        when x"20DB" => data_out<= x"A9";
        when x"20DC" => data_out<= x"FF";
        when x"20DD" => data_out<= x"20";
        when x"20DE" => data_out<= x"65";
        when x"20DF" => data_out<= x"9F";
        when x"20E0" => data_out<= x"A9";
        when x"20E1" => data_out<= x"FF";
        when x"20E2" => data_out<= x"20";
        when x"20E3" => data_out<= x"65";
        when x"20E4" => data_out<= x"9F";
        when x"20E5" => data_out<= x"A9";
        when x"20E6" => data_out<= x"FF";
        when x"20E7" => data_out<= x"20";
        when x"20E8" => data_out<= x"65";
        when x"20E9" => data_out<= x"9F";
        when x"20EA" => data_out<= x"A0";
        when x"20EB" => data_out<= x"00";
        when x"20EC" => data_out<= x"B1";
        when x"20ED" => data_out<= x"0C";
        when x"20EE" => data_out<= x"29";
        when x"20EF" => data_out<= x"40";
        when x"20F0" => data_out<= x"D0";
        when x"20F1" => data_out<= x"05";
        when x"20F2" => data_out<= x"A9";
        when x"20F3" => data_out<= x"01";
        when x"20F4" => data_out<= x"8D";
        when x"20F5" => data_out<= x"04";
        when x"20F6" => data_out<= x"02";
        when x"20F7" => data_out<= x"20";
        when x"20F8" => data_out<= x"05";
        when x"20F9" => data_out<= x"AF";
        when x"20FA" => data_out<= x"20";
        when x"20FB" => data_out<= x"7C";
        when x"20FC" => data_out<= x"A2";
        when x"20FD" => data_out<= x"A9";
        when x"20FE" => data_out<= x"FF";
        when x"20FF" => data_out<= x"20";
        when x"2100" => data_out<= x"65";
        when x"2101" => data_out<= x"9F";
        when x"2102" => data_out<= x"A9";
        when x"2103" => data_out<= x"01";
        when x"2104" => data_out<= x"8D";
        when x"2105" => data_out<= x"05";
        when x"2106" => data_out<= x"02";
        when x"2107" => data_out<= x"A2";
        when x"2108" => data_out<= x"00";
        when x"2109" => data_out<= x"8A";
        when x"210A" => data_out<= x"4C";
        when x"210B" => data_out<= x"27";
        when x"210C" => data_out<= x"AF";
        when x"210D" => data_out<= x"20";
        when x"210E" => data_out<= x"7B";
        when x"210F" => data_out<= x"B0";
        when x"2110" => data_out<= x"20";
        when x"2111" => data_out<= x"80";
        when x"2112" => data_out<= x"AE";
        when x"2113" => data_out<= x"AD";
        when x"2114" => data_out<= x"04";
        when x"2115" => data_out<= x"02";
        when x"2116" => data_out<= x"C9";
        when x"2117" => data_out<= x"02";
        when x"2118" => data_out<= x"F0";
        when x"2119" => data_out<= x"16";
        when x"211A" => data_out<= x"A0";
        when x"211B" => data_out<= x"08";
        when x"211C" => data_out<= x"20";
        when x"211D" => data_out<= x"58";
        when x"211E" => data_out<= x"AF";
        when x"211F" => data_out<= x"A4";
        when x"2120" => data_out<= x"0E";
        when x"2121" => data_out<= x"84";
        when x"2122" => data_out<= x"0F";
        when x"2123" => data_out<= x"86";
        when x"2124" => data_out<= x"0E";
        when x"2125" => data_out<= x"AA";
        when x"2126" => data_out<= x"A9";
        when x"2127" => data_out<= x"00";
        when x"2128" => data_out<= x"20";
        when x"2129" => data_out<= x"3A";
        when x"212A" => data_out<= x"AE";
        when x"212B" => data_out<= x"A0";
        when x"212C" => data_out<= x"05";
        when x"212D" => data_out<= x"20";
        when x"212E" => data_out<= x"EB";
        when x"212F" => data_out<= x"B0";
        when x"2130" => data_out<= x"20";
        when x"2131" => data_out<= x"77";
        when x"2132" => data_out<= x"A2";
        when x"2133" => data_out<= x"A9";
        when x"2134" => data_out<= x"51";
        when x"2135" => data_out<= x"20";
        when x"2136" => data_out<= x"65";
        when x"2137" => data_out<= x"B0";
        when x"2138" => data_out<= x"A0";
        when x"2139" => data_out<= x"09";
        when x"213A" => data_out<= x"20";
        when x"213B" => data_out<= x"58";
        when x"213C" => data_out<= x"AF";
        when x"213D" => data_out<= x"20";
        when x"213E" => data_out<= x"7E";
        when x"213F" => data_out<= x"AF";
        when x"2140" => data_out<= x"A9";
        when x"2141" => data_out<= x"FF";
        when x"2142" => data_out<= x"20";
        when x"2143" => data_out<= x"7F";
        when x"2144" => data_out<= x"A2";
        when x"2145" => data_out<= x"A0";
        when x"2146" => data_out<= x"02";
        when x"2147" => data_out<= x"91";
        when x"2148" => data_out<= x"0C";
        when x"2149" => data_out<= x"A2";
        when x"214A" => data_out<= x"00";
        when x"214B" => data_out<= x"B1";
        when x"214C" => data_out<= x"0C";
        when x"214D" => data_out<= x"F0";
        when x"214E" => data_out<= x"0A";
        when x"214F" => data_out<= x"20";
        when x"2150" => data_out<= x"7C";
        when x"2151" => data_out<= x"A2";
        when x"2152" => data_out<= x"A2";
        when x"2153" => data_out<= x"00";
        when x"2154" => data_out<= x"A9";
        when x"2155" => data_out<= x"02";
        when x"2156" => data_out<= x"4C";
        when x"2157" => data_out<= x"B0";
        when x"2158" => data_out<= x"A1";
        when x"2159" => data_out<= x"20";
        when x"215A" => data_out<= x"C3";
        when x"215B" => data_out<= x"B0";
        when x"215C" => data_out<= x"A0";
        when x"215D" => data_out<= x"01";
        when x"215E" => data_out<= x"B1";
        when x"215F" => data_out<= x"0C";
        when x"2160" => data_out<= x"C9";
        when x"2161" => data_out<= x"13";
        when x"2162" => data_out<= x"D0";
        when x"2163" => data_out<= x"05";
        when x"2164" => data_out<= x"88";
        when x"2165" => data_out<= x"B1";
        when x"2166" => data_out<= x"0C";
        when x"2167" => data_out<= x"C9";
        when x"2168" => data_out<= x"88";
        when x"2169" => data_out<= x"B0";
        when x"216A" => data_out<= x"16";
        when x"216B" => data_out<= x"A9";
        when x"216C" => data_out<= x"FF";
        when x"216D" => data_out<= x"20";
        when x"216E" => data_out<= x"65";
        when x"216F" => data_out<= x"9F";
        when x"2170" => data_out<= x"A0";
        when x"2171" => data_out<= x"02";
        when x"2172" => data_out<= x"91";
        when x"2173" => data_out<= x"0C";
        when x"2174" => data_out<= x"C9";
        when x"2175" => data_out<= x"FE";
        when x"2176" => data_out<= x"F0";
        when x"2177" => data_out<= x"0B";
        when x"2178" => data_out<= x"20";
        when x"2179" => data_out<= x"4D";
        when x"217A" => data_out<= x"AF";
        when x"217B" => data_out<= x"20";
        when x"217C" => data_out<= x"E2";
        when x"217D" => data_out<= x"AE";
        when x"217E" => data_out<= x"4C";
        when x"217F" => data_out<= x"59";
        when x"2180" => data_out<= x"A1";
        when x"2181" => data_out<= x"A0";
        when x"2182" => data_out<= x"02";
        when x"2183" => data_out<= x"B1";
        when x"2184" => data_out<= x"0C";
        when x"2185" => data_out<= x"C9";
        when x"2186" => data_out<= x"FE";
        when x"2187" => data_out<= x"F0";
        when x"2188" => data_out<= x"0A";
        when x"2189" => data_out<= x"20";
        when x"218A" => data_out<= x"7C";
        when x"218B" => data_out<= x"A2";
        when x"218C" => data_out<= x"A2";
        when x"218D" => data_out<= x"00";
        when x"218E" => data_out<= x"A9";
        when x"218F" => data_out<= x"01";
        when x"2190" => data_out<= x"4C";
        when x"2191" => data_out<= x"B0";
        when x"2192" => data_out<= x"A1";
        when x"2193" => data_out<= x"A0";
        when x"2194" => data_out<= x"04";
        when x"2195" => data_out<= x"20";
        when x"2196" => data_out<= x"4F";
        when x"2197" => data_out<= x"AF";
        when x"2198" => data_out<= x"20";
        when x"2199" => data_out<= x"18";
        when x"219A" => data_out<= x"A3";
        when x"219B" => data_out<= x"A9";
        when x"219C" => data_out<= x"FF";
        when x"219D" => data_out<= x"20";
        when x"219E" => data_out<= x"65";
        when x"219F" => data_out<= x"9F";
        when x"21A0" => data_out<= x"A9";
        when x"21A1" => data_out<= x"FF";
        when x"21A2" => data_out<= x"20";
        when x"21A3" => data_out<= x"65";
        when x"21A4" => data_out<= x"9F";
        when x"21A5" => data_out<= x"20";
        when x"21A6" => data_out<= x"7C";
        when x"21A7" => data_out<= x"A2";
        when x"21A8" => data_out<= x"A9";
        when x"21A9" => data_out<= x"FF";
        when x"21AA" => data_out<= x"20";
        when x"21AB" => data_out<= x"65";
        when x"21AC" => data_out<= x"9F";
        when x"21AD" => data_out<= x"A2";
        when x"21AE" => data_out<= x"00";
        when x"21AF" => data_out<= x"8A";
        when x"21B0" => data_out<= x"A0";
        when x"21B1" => data_out<= x"09";
        when x"21B2" => data_out<= x"4C";
        when x"21B3" => data_out<= x"14";
        when x"21B4" => data_out<= x"AE";
        when x"21B5" => data_out<= x"20";
        when x"21B6" => data_out<= x"7B";
        when x"21B7" => data_out<= x"B0";
        when x"21B8" => data_out<= x"20";
        when x"21B9" => data_out<= x"80";
        when x"21BA" => data_out<= x"AE";
        when x"21BB" => data_out<= x"AD";
        when x"21BC" => data_out<= x"04";
        when x"21BD" => data_out<= x"02";
        when x"21BE" => data_out<= x"C9";
        when x"21BF" => data_out<= x"02";
        when x"21C0" => data_out<= x"F0";
        when x"21C1" => data_out<= x"16";
        when x"21C2" => data_out<= x"A0";
        when x"21C3" => data_out<= x"08";
        when x"21C4" => data_out<= x"20";
        when x"21C5" => data_out<= x"58";
        when x"21C6" => data_out<= x"AF";
        when x"21C7" => data_out<= x"A4";
        when x"21C8" => data_out<= x"0E";
        when x"21C9" => data_out<= x"84";
        when x"21CA" => data_out<= x"0F";
        when x"21CB" => data_out<= x"86";
        when x"21CC" => data_out<= x"0E";
        when x"21CD" => data_out<= x"AA";
        when x"21CE" => data_out<= x"A9";
        when x"21CF" => data_out<= x"00";
        when x"21D0" => data_out<= x"20";
        when x"21D1" => data_out<= x"3A";
        when x"21D2" => data_out<= x"AE";
        when x"21D3" => data_out<= x"A0";
        when x"21D4" => data_out<= x"05";
        when x"21D5" => data_out<= x"20";
        when x"21D6" => data_out<= x"EB";
        when x"21D7" => data_out<= x"B0";
        when x"21D8" => data_out<= x"20";
        when x"21D9" => data_out<= x"77";
        when x"21DA" => data_out<= x"A2";
        when x"21DB" => data_out<= x"A9";
        when x"21DC" => data_out<= x"58";
        when x"21DD" => data_out<= x"20";
        when x"21DE" => data_out<= x"65";
        when x"21DF" => data_out<= x"B0";
        when x"21E0" => data_out<= x"A0";
        when x"21E1" => data_out<= x"09";
        when x"21E2" => data_out<= x"20";
        when x"21E3" => data_out<= x"58";
        when x"21E4" => data_out<= x"AF";
        when x"21E5" => data_out<= x"20";
        when x"21E6" => data_out<= x"7E";
        when x"21E7" => data_out<= x"AF";
        when x"21E8" => data_out<= x"A9";
        when x"21E9" => data_out<= x"FF";
        when x"21EA" => data_out<= x"20";
        when x"21EB" => data_out<= x"7F";
        when x"21EC" => data_out<= x"A2";
        when x"21ED" => data_out<= x"A0";
        when x"21EE" => data_out<= x"02";
        when x"21EF" => data_out<= x"91";
        when x"21F0" => data_out<= x"0C";
        when x"21F1" => data_out<= x"B1";
        when x"21F2" => data_out<= x"0C";
        when x"21F3" => data_out<= x"F0";
        when x"21F4" => data_out<= x"0A";
        when x"21F5" => data_out<= x"20";
        when x"21F6" => data_out<= x"7C";
        when x"21F7" => data_out<= x"A2";
        when x"21F8" => data_out<= x"A2";
        when x"21F9" => data_out<= x"00";
        when x"21FA" => data_out<= x"A9";
        when x"21FB" => data_out<= x"02";
        when x"21FC" => data_out<= x"4C";
        when x"21FD" => data_out<= x"66";
        when x"21FE" => data_out<= x"A2";
        when x"21FF" => data_out<= x"A9";
        when x"2200" => data_out<= x"FF";
        when x"2201" => data_out<= x"20";
        when x"2202" => data_out<= x"65";
        when x"2203" => data_out<= x"9F";
        when x"2204" => data_out<= x"A9";
        when x"2205" => data_out<= x"FE";
        when x"2206" => data_out<= x"20";
        when x"2207" => data_out<= x"65";
        when x"2208" => data_out<= x"9F";
        when x"2209" => data_out<= x"A0";
        when x"220A" => data_out<= x"04";
        when x"220B" => data_out<= x"20";
        when x"220C" => data_out<= x"4F";
        when x"220D" => data_out<= x"AF";
        when x"220E" => data_out<= x"20";
        when x"220F" => data_out<= x"41";
        when x"2210" => data_out<= x"A3";
        when x"2211" => data_out<= x"A9";
        when x"2212" => data_out<= x"FF";
        when x"2213" => data_out<= x"20";
        when x"2214" => data_out<= x"65";
        when x"2215" => data_out<= x"9F";
        when x"2216" => data_out<= x"A9";
        when x"2217" => data_out<= x"FF";
        when x"2218" => data_out<= x"20";
        when x"2219" => data_out<= x"65";
        when x"221A" => data_out<= x"9F";
        when x"221B" => data_out<= x"A9";
        when x"221C" => data_out<= x"FF";
        when x"221D" => data_out<= x"20";
        when x"221E" => data_out<= x"65";
        when x"221F" => data_out<= x"9F";
        when x"2220" => data_out<= x"A0";
        when x"2221" => data_out<= x"02";
        when x"2222" => data_out<= x"91";
        when x"2223" => data_out<= x"0C";
        when x"2224" => data_out<= x"A2";
        when x"2225" => data_out<= x"00";
        when x"2226" => data_out<= x"29";
        when x"2227" => data_out<= x"1F";
        when x"2228" => data_out<= x"C9";
        when x"2229" => data_out<= x"05";
        when x"222A" => data_out<= x"F0";
        when x"222B" => data_out<= x"0A";
        when x"222C" => data_out<= x"20";
        when x"222D" => data_out<= x"7C";
        when x"222E" => data_out<= x"A2";
        when x"222F" => data_out<= x"A2";
        when x"2230" => data_out<= x"00";
        when x"2231" => data_out<= x"A9";
        when x"2232" => data_out<= x"05";
        when x"2233" => data_out<= x"4C";
        when x"2234" => data_out<= x"66";
        when x"2235" => data_out<= x"A2";
        when x"2236" => data_out<= x"8A";
        when x"2237" => data_out<= x"20";
        when x"2238" => data_out<= x"C3";
        when x"2239" => data_out<= x"B0";
        when x"223A" => data_out<= x"A0";
        when x"223B" => data_out<= x"01";
        when x"223C" => data_out<= x"B1";
        when x"223D" => data_out<= x"0C";
        when x"223E" => data_out<= x"C9";
        when x"223F" => data_out<= x"27";
        when x"2240" => data_out<= x"D0";
        when x"2241" => data_out<= x"05";
        when x"2242" => data_out<= x"88";
        when x"2243" => data_out<= x"B1";
        when x"2244" => data_out<= x"0C";
        when x"2245" => data_out<= x"C9";
        when x"2246" => data_out<= x"10";
        when x"2247" => data_out<= x"B0";
        when x"2248" => data_out<= x"12";
        when x"2249" => data_out<= x"A9";
        when x"224A" => data_out<= x"FF";
        when x"224B" => data_out<= x"20";
        when x"224C" => data_out<= x"65";
        when x"224D" => data_out<= x"9F";
        when x"224E" => data_out<= x"C9";
        when x"224F" => data_out<= x"00";
        when x"2250" => data_out<= x"D0";
        when x"2251" => data_out<= x"09";
        when x"2252" => data_out<= x"20";
        when x"2253" => data_out<= x"4D";
        when x"2254" => data_out<= x"AF";
        when x"2255" => data_out<= x"20";
        when x"2256" => data_out<= x"E2";
        when x"2257" => data_out<= x"AE";
        when x"2258" => data_out<= x"4C";
        when x"2259" => data_out<= x"37";
        when x"225A" => data_out<= x"A2";
        when x"225B" => data_out<= x"20";
        when x"225C" => data_out<= x"7C";
        when x"225D" => data_out<= x"A2";
        when x"225E" => data_out<= x"A9";
        when x"225F" => data_out<= x"FF";
        when x"2260" => data_out<= x"20";
        when x"2261" => data_out<= x"65";
        when x"2262" => data_out<= x"9F";
        when x"2263" => data_out<= x"A2";
        when x"2264" => data_out<= x"00";
        when x"2265" => data_out<= x"8A";
        when x"2266" => data_out<= x"A0";
        when x"2267" => data_out<= x"09";
        when x"2268" => data_out<= x"4C";
        when x"2269" => data_out<= x"14";
        when x"226A" => data_out<= x"AE";
        when x"226B" => data_out<= x"A2";
        when x"226C" => data_out<= x"00";
        when x"226D" => data_out<= x"AD";
        when x"226E" => data_out<= x"05";
        when x"226F" => data_out<= x"02";
        when x"2270" => data_out<= x"60";
        when x"2271" => data_out<= x"A2";
        when x"2272" => data_out<= x"00";
        when x"2273" => data_out<= x"AD";
        when x"2274" => data_out<= x"04";
        when x"2275" => data_out<= x"02";
        when x"2276" => data_out<= x"60";
        when x"2277" => data_out<= x"A9";
        when x"2278" => data_out<= x"01";
        when x"2279" => data_out<= x"4C";
        when x"227A" => data_out<= x"56";
        when x"227B" => data_out<= x"9F";
        when x"227C" => data_out<= x"4C";
        when x"227D" => data_out<= x"5F";
        when x"227E" => data_out<= x"9F";
        when x"227F" => data_out<= x"20";
        when x"2280" => data_out<= x"65";
        when x"2281" => data_out<= x"B0";
        when x"2282" => data_out<= x"20";
        when x"2283" => data_out<= x"73";
        when x"2284" => data_out<= x"AE";
        when x"2285" => data_out<= x"A9";
        when x"2286" => data_out<= x"FF";
        when x"2287" => data_out<= x"20";
        when x"2288" => data_out<= x"65";
        when x"2289" => data_out<= x"9F";
        when x"228A" => data_out<= x"A0";
        when x"228B" => data_out<= x"07";
        when x"228C" => data_out<= x"B1";
        when x"228D" => data_out<= x"0C";
        when x"228E" => data_out<= x"20";
        when x"228F" => data_out<= x"65";
        when x"2290" => data_out<= x"9F";
        when x"2291" => data_out<= x"A0";
        when x"2292" => data_out<= x"06";
        when x"2293" => data_out<= x"20";
        when x"2294" => data_out<= x"58";
        when x"2295" => data_out<= x"AF";
        when x"2296" => data_out<= x"A5";
        when x"2297" => data_out<= x"0F";
        when x"2298" => data_out<= x"20";
        when x"2299" => data_out<= x"65";
        when x"229A" => data_out<= x"9F";
        when x"229B" => data_out<= x"A0";
        when x"229C" => data_out<= x"06";
        when x"229D" => data_out<= x"20";
        when x"229E" => data_out<= x"58";
        when x"229F" => data_out<= x"AF";
        when x"22A0" => data_out<= x"A5";
        when x"22A1" => data_out<= x"0E";
        when x"22A2" => data_out<= x"20";
        when x"22A3" => data_out<= x"65";
        when x"22A4" => data_out<= x"9F";
        when x"22A5" => data_out<= x"A0";
        when x"22A6" => data_out<= x"06";
        when x"22A7" => data_out<= x"20";
        when x"22A8" => data_out<= x"58";
        when x"22A9" => data_out<= x"AF";
        when x"22AA" => data_out<= x"8A";
        when x"22AB" => data_out<= x"20";
        when x"22AC" => data_out<= x"65";
        when x"22AD" => data_out<= x"9F";
        when x"22AE" => data_out<= x"A0";
        when x"22AF" => data_out<= x"06";
        when x"22B0" => data_out<= x"20";
        when x"22B1" => data_out<= x"58";
        when x"22B2" => data_out<= x"AF";
        when x"22B3" => data_out<= x"20";
        when x"22B4" => data_out<= x"65";
        when x"22B5" => data_out<= x"9F";
        when x"22B6" => data_out<= x"A0";
        when x"22B7" => data_out<= x"02";
        when x"22B8" => data_out<= x"B1";
        when x"22B9" => data_out<= x"0C";
        when x"22BA" => data_out<= x"20";
        when x"22BB" => data_out<= x"65";
        when x"22BC" => data_out<= x"9F";
        when x"22BD" => data_out<= x"A9";
        when x"22BE" => data_out<= x"00";
        when x"22BF" => data_out<= x"A8";
        when x"22C0" => data_out<= x"91";
        when x"22C1" => data_out<= x"0C";
        when x"22C2" => data_out<= x"AA";
        when x"22C3" => data_out<= x"B1";
        when x"22C4" => data_out<= x"0C";
        when x"22C5" => data_out<= x"C9";
        when x"22C6" => data_out<= x"0A";
        when x"22C7" => data_out<= x"B0";
        when x"22C8" => data_out<= x"21";
        when x"22C9" => data_out<= x"A9";
        when x"22CA" => data_out<= x"FF";
        when x"22CB" => data_out<= x"20";
        when x"22CC" => data_out<= x"65";
        when x"22CD" => data_out<= x"9F";
        when x"22CE" => data_out<= x"A0";
        when x"22CF" => data_out<= x"01";
        when x"22D0" => data_out<= x"91";
        when x"22D1" => data_out<= x"0C";
        when x"22D2" => data_out<= x"C9";
        when x"22D3" => data_out<= x"FF";
        when x"22D4" => data_out<= x"F0";
        when x"22D5" => data_out<= x"07";
        when x"22D6" => data_out<= x"A2";
        when x"22D7" => data_out<= x"00";
        when x"22D8" => data_out<= x"B1";
        when x"22D9" => data_out<= x"0C";
        when x"22DA" => data_out<= x"4C";
        when x"22DB" => data_out<= x"3B";
        when x"22DC" => data_out<= x"AF";
        when x"22DD" => data_out<= x"88";
        when x"22DE" => data_out<= x"A2";
        when x"22DF" => data_out<= x"00";
        when x"22E0" => data_out<= x"B1";
        when x"22E1" => data_out<= x"0C";
        when x"22E2" => data_out<= x"18";
        when x"22E3" => data_out<= x"69";
        when x"22E4" => data_out<= x"01";
        when x"22E5" => data_out<= x"91";
        when x"22E6" => data_out<= x"0C";
        when x"22E7" => data_out<= x"4C";
        when x"22E8" => data_out<= x"C3";
        when x"22E9" => data_out<= x"A2";
        when x"22EA" => data_out<= x"A9";
        when x"22EB" => data_out<= x"FF";
        when x"22EC" => data_out<= x"4C";
        when x"22ED" => data_out<= x"3B";
        when x"22EE" => data_out<= x"AF";
        when x"22EF" => data_out<= x"20";
        when x"22F0" => data_out<= x"7E";
        when x"22F1" => data_out<= x"AF";
        when x"22F2" => data_out<= x"A9";
        when x"22F3" => data_out<= x"77";
        when x"22F4" => data_out<= x"20";
        when x"22F5" => data_out<= x"65";
        when x"22F6" => data_out<= x"B0";
        when x"22F7" => data_out<= x"A2";
        when x"22F8" => data_out<= x"00";
        when x"22F9" => data_out<= x"20";
        when x"22FA" => data_out<= x"75";
        when x"22FB" => data_out<= x"AF";
        when x"22FC" => data_out<= x"A9";
        when x"22FD" => data_out<= x"65";
        when x"22FE" => data_out<= x"20";
        when x"22FF" => data_out<= x"7F";
        when x"2300" => data_out<= x"A2";
        when x"2301" => data_out<= x"A0";
        when x"2302" => data_out<= x"04";
        when x"2303" => data_out<= x"B1";
        when x"2304" => data_out<= x"0C";
        when x"2305" => data_out<= x"20";
        when x"2306" => data_out<= x"65";
        when x"2307" => data_out<= x"B0";
        when x"2308" => data_out<= x"A0";
        when x"2309" => data_out<= x"04";
        when x"230A" => data_out<= x"20";
        when x"230B" => data_out<= x"58";
        when x"230C" => data_out<= x"AF";
        when x"230D" => data_out<= x"20";
        when x"230E" => data_out<= x"7E";
        when x"230F" => data_out<= x"AF";
        when x"2310" => data_out<= x"A9";
        when x"2311" => data_out<= x"FF";
        when x"2312" => data_out<= x"20";
        when x"2313" => data_out<= x"7F";
        when x"2314" => data_out<= x"A2";
        when x"2315" => data_out<= x"4C";
        when x"2316" => data_out<= x"2C";
        when x"2317" => data_out<= x"AF";
        when x"2318" => data_out<= x"85";
        when x"2319" => data_out<= x"14";
        when x"231A" => data_out<= x"86";
        when x"231B" => data_out<= x"15";
        when x"231C" => data_out<= x"A2";
        when x"231D" => data_out<= x"02";
        when x"231E" => data_out<= x"A0";
        when x"231F" => data_out<= x"00";
        when x"2320" => data_out<= x"AD";
        when x"2321" => data_out<= x"42";
        when x"2322" => data_out<= x"C0";
        when x"2323" => data_out<= x"29";
        when x"2324" => data_out<= x"20";
        when x"2325" => data_out<= x"F0";
        when x"2326" => data_out<= x"F9";
        when x"2327" => data_out<= x"A9";
        when x"2328" => data_out<= x"FF";
        when x"2329" => data_out<= x"8D";
        when x"232A" => data_out<= x"41";
        when x"232B" => data_out<= x"C0";
        when x"232C" => data_out<= x"AD";
        when x"232D" => data_out<= x"42";
        when x"232E" => data_out<= x"C0";
        when x"232F" => data_out<= x"29";
        when x"2330" => data_out<= x"40";
        when x"2331" => data_out<= x"F0";
        when x"2332" => data_out<= x"F9";
        when x"2333" => data_out<= x"AD";
        when x"2334" => data_out<= x"40";
        when x"2335" => data_out<= x"C0";
        when x"2336" => data_out<= x"91";
        when x"2337" => data_out<= x"14";
        when x"2338" => data_out<= x"C8";
        when x"2339" => data_out<= x"D0";
        when x"233A" => data_out<= x"E5";
        when x"233B" => data_out<= x"E6";
        when x"233C" => data_out<= x"15";
        when x"233D" => data_out<= x"CA";
        when x"233E" => data_out<= x"D0";
        when x"233F" => data_out<= x"E0";
        when x"2340" => data_out<= x"60";
        when x"2341" => data_out<= x"85";
        when x"2342" => data_out<= x"14";
        when x"2343" => data_out<= x"86";
        when x"2344" => data_out<= x"15";
        when x"2345" => data_out<= x"A2";
        when x"2346" => data_out<= x"02";
        when x"2347" => data_out<= x"A0";
        when x"2348" => data_out<= x"00";
        when x"2349" => data_out<= x"AD";
        when x"234A" => data_out<= x"42";
        when x"234B" => data_out<= x"C0";
        when x"234C" => data_out<= x"29";
        when x"234D" => data_out<= x"20";
        when x"234E" => data_out<= x"F0";
        when x"234F" => data_out<= x"F9";
        when x"2350" => data_out<= x"B1";
        when x"2351" => data_out<= x"14";
        when x"2352" => data_out<= x"8D";
        when x"2353" => data_out<= x"41";
        when x"2354" => data_out<= x"C0";
        when x"2355" => data_out<= x"AD";
        when x"2356" => data_out<= x"42";
        when x"2357" => data_out<= x"C0";
        when x"2358" => data_out<= x"29";
        when x"2359" => data_out<= x"40";
        when x"235A" => data_out<= x"F0";
        when x"235B" => data_out<= x"F9";
        when x"235C" => data_out<= x"AD";
        when x"235D" => data_out<= x"40";
        when x"235E" => data_out<= x"C0";
        when x"235F" => data_out<= x"C8";
        when x"2360" => data_out<= x"D0";
        when x"2361" => data_out<= x"E7";
        when x"2362" => data_out<= x"E6";
        when x"2363" => data_out<= x"15";
        when x"2364" => data_out<= x"CA";
        when x"2365" => data_out<= x"D0";
        when x"2366" => data_out<= x"E2";
        when x"2367" => data_out<= x"60";
        when x"2368" => data_out<= x"A9";
        when x"2369" => data_out<= x"00";
        when x"236A" => data_out<= x"8D";
        when x"236B" => data_out<= x"47";
        when x"236C" => data_out<= x"02";
        when x"236D" => data_out<= x"20";
        when x"236E" => data_out<= x"BF";
        when x"236F" => data_out<= x"9F";
        when x"2370" => data_out<= x"AA";
        when x"2371" => data_out<= x"F0";
        when x"2372" => data_out<= x"05";
        when x"2373" => data_out<= x"A2";
        when x"2374" => data_out<= x"00";
        when x"2375" => data_out<= x"A9";
        when x"2376" => data_out<= x"01";
        when x"2377" => data_out<= x"60";
        when x"2378" => data_out<= x"20";
        when x"2379" => data_out<= x"75";
        when x"237A" => data_out<= x"AF";
        when x"237B" => data_out<= x"A9";
        when x"237C" => data_out<= x"54";
        when x"237D" => data_out<= x"A2";
        when x"237E" => data_out<= x"02";
        when x"237F" => data_out<= x"20";
        when x"2380" => data_out<= x"0D";
        when x"2381" => data_out<= x"A1";
        when x"2382" => data_out<= x"AA";
        when x"2383" => data_out<= x"F0";
        when x"2384" => data_out<= x"05";
        when x"2385" => data_out<= x"A2";
        when x"2386" => data_out<= x"00";
        when x"2387" => data_out<= x"A9";
        when x"2388" => data_out<= x"01";
        when x"2389" => data_out<= x"60";
        when x"238A" => data_out<= x"AD";
        when x"238B" => data_out<= x"54";
        when x"238C" => data_out<= x"02";
        when x"238D" => data_out<= x"C9";
        when x"238E" => data_out<= x"46";
        when x"238F" => data_out<= x"D0";
        when x"2390" => data_out<= x"09";
        when x"2391" => data_out<= x"AD";
        when x"2392" => data_out<= x"55";
        when x"2393" => data_out<= x"02";
        when x"2394" => data_out<= x"C9";
        when x"2395" => data_out<= x"4D";
        when x"2396" => data_out<= x"D0";
        when x"2397" => data_out<= x"02";
        when x"2398" => data_out<= x"8A";
        when x"2399" => data_out<= x"60";
        when x"239A" => data_out<= x"A9";
        when x"239B" => data_out<= x"02";
        when x"239C" => data_out<= x"60";
        when x"239D" => data_out<= x"A9";
        when x"239E" => data_out<= x"00";
        when x"239F" => data_out<= x"8D";
        when x"23A0" => data_out<= x"47";
        when x"23A1" => data_out<= x"02";
        when x"23A2" => data_out<= x"20";
        when x"23A3" => data_out<= x"BF";
        when x"23A4" => data_out<= x"9F";
        when x"23A5" => data_out<= x"AA";
        when x"23A6" => data_out<= x"F0";
        when x"23A7" => data_out<= x"05";
        when x"23A8" => data_out<= x"A2";
        when x"23A9" => data_out<= x"00";
        when x"23AA" => data_out<= x"A9";
        when x"23AB" => data_out<= x"01";
        when x"23AC" => data_out<= x"60";
        when x"23AD" => data_out<= x"A9";
        when x"23AE" => data_out<= x"54";
        when x"23AF" => data_out<= x"A2";
        when x"23B0" => data_out<= x"02";
        when x"23B1" => data_out<= x"20";
        when x"23B2" => data_out<= x"7B";
        when x"23B3" => data_out<= x"B0";
        when x"23B4" => data_out<= x"A2";
        when x"23B5" => data_out<= x"02";
        when x"23B6" => data_out<= x"A9";
        when x"23B7" => data_out<= x"00";
        when x"23B8" => data_out<= x"20";
        when x"23B9" => data_out<= x"D2";
        when x"23BA" => data_out<= x"AF";
        when x"23BB" => data_out<= x"A9";
        when x"23BC" => data_out<= x"46";
        when x"23BD" => data_out<= x"8D";
        when x"23BE" => data_out<= x"54";
        when x"23BF" => data_out<= x"02";
        when x"23C0" => data_out<= x"A9";
        when x"23C1" => data_out<= x"4D";
        when x"23C2" => data_out<= x"8D";
        when x"23C3" => data_out<= x"55";
        when x"23C4" => data_out<= x"02";
        when x"23C5" => data_out<= x"A9";
        when x"23C6" => data_out<= x"01";
        when x"23C7" => data_out<= x"8D";
        when x"23C8" => data_out<= x"5A";
        when x"23C9" => data_out<= x"02";
        when x"23CA" => data_out<= x"A9";
        when x"23CB" => data_out<= x"00";
        when x"23CC" => data_out<= x"8D";
        when x"23CD" => data_out<= x"5B";
        when x"23CE" => data_out<= x"02";
        when x"23CF" => data_out<= x"20";
        when x"23D0" => data_out<= x"37";
        when x"23D1" => data_out<= x"AB";
        when x"23D2" => data_out<= x"86";
        when x"23D3" => data_out<= x"1C";
        when x"23D4" => data_out<= x"05";
        when x"23D5" => data_out<= x"1C";
        when x"23D6" => data_out<= x"F0";
        when x"23D7" => data_out<= x"05";
        when x"23D8" => data_out<= x"A2";
        when x"23D9" => data_out<= x"00";
        when x"23DA" => data_out<= x"A9";
        when x"23DB" => data_out<= x"01";
        when x"23DC" => data_out<= x"60";
        when x"23DD" => data_out<= x"A2";
        when x"23DE" => data_out<= x"00";
        when x"23DF" => data_out<= x"60";
        when x"23E0" => data_out<= x"20";
        when x"23E1" => data_out<= x"7B";
        when x"23E2" => data_out<= x"B0";
        when x"23E3" => data_out<= x"20";
        when x"23E4" => data_out<= x"80";
        when x"23E5" => data_out<= x"AE";
        when x"23E6" => data_out<= x"20";
        when x"23E7" => data_out<= x"B9";
        when x"23E8" => data_out<= x"A9";
        when x"23E9" => data_out<= x"A9";
        when x"23EA" => data_out<= x"00";
        when x"23EB" => data_out<= x"A0";
        when x"23EC" => data_out<= x"02";
        when x"23ED" => data_out<= x"91";
        when x"23EE" => data_out<= x"0C";
        when x"23EF" => data_out<= x"AA";
        when x"23F0" => data_out<= x"B1";
        when x"23F1" => data_out<= x"0C";
        when x"23F2" => data_out<= x"C9";
        when x"23F3" => data_out<= x"10";
        when x"23F4" => data_out<= x"90";
        when x"23F5" => data_out<= x"03";
        when x"23F6" => data_out<= x"4C";
        when x"23F7" => data_out<= x"B7";
        when x"23F8" => data_out<= x"A4";
        when x"23F9" => data_out<= x"20";
        when x"23FA" => data_out<= x"29";
        when x"23FB" => data_out<= x"AE";
        when x"23FC" => data_out<= x"20";
        when x"23FD" => data_out<= x"21";
        when x"23FE" => data_out<= x"AE";
        when x"23FF" => data_out<= x"18";
        when x"2400" => data_out<= x"69";
        when x"2401" => data_out<= x"64";
        when x"2402" => data_out<= x"A8";
        when x"2403" => data_out<= x"8A";
        when x"2404" => data_out<= x"69";
        when x"2405" => data_out<= x"02";
        when x"2406" => data_out<= x"AA";
        when x"2407" => data_out<= x"98";
        when x"2408" => data_out<= x"20";
        when x"2409" => data_out<= x"C3";
        when x"240A" => data_out<= x"B0";
        when x"240B" => data_out<= x"85";
        when x"240C" => data_out<= x"14";
        when x"240D" => data_out<= x"86";
        when x"240E" => data_out<= x"15";
        when x"240F" => data_out<= x"A0";
        when x"2410" => data_out<= x"00";
        when x"2411" => data_out<= x"B1";
        when x"2412" => data_out<= x"14";
        when x"2413" => data_out<= x"D0";
        when x"2414" => data_out<= x"03";
        when x"2415" => data_out<= x"4C";
        when x"2416" => data_out<= x"AA";
        when x"2417" => data_out<= x"A4";
        when x"2418" => data_out<= x"20";
        when x"2419" => data_out<= x"91";
        when x"241A" => data_out<= x"B0";
        when x"241B" => data_out<= x"A0";
        when x"241C" => data_out<= x"06";
        when x"241D" => data_out<= x"20";
        when x"241E" => data_out<= x"4F";
        when x"241F" => data_out<= x"AF";
        when x"2420" => data_out<= x"20";
        when x"2421" => data_out<= x"43";
        when x"2422" => data_out<= x"AB";
        when x"2423" => data_out<= x"AA";
        when x"2424" => data_out<= x"D0";
        when x"2425" => data_out<= x"03";
        when x"2426" => data_out<= x"4C";
        when x"2427" => data_out<= x"AA";
        when x"2428" => data_out<= x"A4";
        when x"2429" => data_out<= x"A0";
        when x"242A" => data_out<= x"02";
        when x"242B" => data_out<= x"B1";
        when x"242C" => data_out<= x"0C";
        when x"242D" => data_out<= x"8D";
        when x"242E" => data_out<= x"49";
        when x"242F" => data_out<= x"02";
        when x"2430" => data_out<= x"20";
        when x"2431" => data_out<= x"4D";
        when x"2432" => data_out<= x"AF";
        when x"2433" => data_out<= x"85";
        when x"2434" => data_out<= x"14";
        when x"2435" => data_out<= x"86";
        when x"2436" => data_out<= x"15";
        when x"2437" => data_out<= x"A0";
        when x"2438" => data_out<= x"0C";
        when x"2439" => data_out<= x"B1";
        when x"243A" => data_out<= x"14";
        when x"243B" => data_out<= x"20";
        when x"243C" => data_out<= x"79";
        when x"243D" => data_out<= x"B0";
        when x"243E" => data_out<= x"A0";
        when x"243F" => data_out<= x"03";
        when x"2440" => data_out<= x"20";
        when x"2441" => data_out<= x"4F";
        when x"2442" => data_out<= x"AF";
        when x"2443" => data_out<= x"85";
        when x"2444" => data_out<= x"14";
        when x"2445" => data_out<= x"86";
        when x"2446" => data_out<= x"15";
        when x"2447" => data_out<= x"A0";
        when x"2448" => data_out<= x"0D";
        when x"2449" => data_out<= x"B1";
        when x"244A" => data_out<= x"14";
        when x"244B" => data_out<= x"AA";
        when x"244C" => data_out<= x"A9";
        when x"244D" => data_out<= x"00";
        when x"244E" => data_out<= x"20";
        when x"244F" => data_out<= x"43";
        when x"2450" => data_out<= x"B0";
        when x"2451" => data_out<= x"8D";
        when x"2452" => data_out<= x"4A";
        when x"2453" => data_out<= x"02";
        when x"2454" => data_out<= x"8E";
        when x"2455" => data_out<= x"4B";
        when x"2456" => data_out<= x"02";
        when x"2457" => data_out<= x"20";
        when x"2458" => data_out<= x"4D";
        when x"2459" => data_out<= x"AF";
        when x"245A" => data_out<= x"85";
        when x"245B" => data_out<= x"14";
        when x"245C" => data_out<= x"86";
        when x"245D" => data_out<= x"15";
        when x"245E" => data_out<= x"A0";
        when x"245F" => data_out<= x"0E";
        when x"2460" => data_out<= x"B1";
        when x"2461" => data_out<= x"14";
        when x"2462" => data_out<= x"20";
        when x"2463" => data_out<= x"79";
        when x"2464" => data_out<= x"B0";
        when x"2465" => data_out<= x"A0";
        when x"2466" => data_out<= x"03";
        when x"2467" => data_out<= x"20";
        when x"2468" => data_out<= x"4F";
        when x"2469" => data_out<= x"AF";
        when x"246A" => data_out<= x"85";
        when x"246B" => data_out<= x"14";
        when x"246C" => data_out<= x"86";
        when x"246D" => data_out<= x"15";
        when x"246E" => data_out<= x"A0";
        when x"246F" => data_out<= x"0F";
        when x"2470" => data_out<= x"B1";
        when x"2471" => data_out<= x"14";
        when x"2472" => data_out<= x"AA";
        when x"2473" => data_out<= x"A9";
        when x"2474" => data_out<= x"00";
        when x"2475" => data_out<= x"20";
        when x"2476" => data_out<= x"43";
        when x"2477" => data_out<= x"B0";
        when x"2478" => data_out<= x"8D";
        when x"2479" => data_out<= x"4C";
        when x"247A" => data_out<= x"02";
        when x"247B" => data_out<= x"8E";
        when x"247C" => data_out<= x"4D";
        when x"247D" => data_out<= x"02";
        when x"247E" => data_out<= x"A9";
        when x"247F" => data_out<= x"00";
        when x"2480" => data_out<= x"8D";
        when x"2481" => data_out<= x"4E";
        when x"2482" => data_out<= x"02";
        when x"2483" => data_out<= x"8D";
        when x"2484" => data_out<= x"4F";
        when x"2485" => data_out<= x"02";
        when x"2486" => data_out<= x"AD";
        when x"2487" => data_out<= x"4B";
        when x"2488" => data_out<= x"02";
        when x"2489" => data_out<= x"8D";
        when x"248A" => data_out<= x"51";
        when x"248B" => data_out<= x"02";
        when x"248C" => data_out<= x"AD";
        when x"248D" => data_out<= x"4A";
        when x"248E" => data_out<= x"02";
        when x"248F" => data_out<= x"8D";
        when x"2490" => data_out<= x"50";
        when x"2491" => data_out<= x"02";
        when x"2492" => data_out<= x"A2";
        when x"2493" => data_out<= x"02";
        when x"2494" => data_out<= x"A9";
        when x"2495" => data_out<= x"00";
        when x"2496" => data_out<= x"8D";
        when x"2497" => data_out<= x"52";
        when x"2498" => data_out<= x"02";
        when x"2499" => data_out<= x"8E";
        when x"249A" => data_out<= x"53";
        when x"249B" => data_out<= x"02";
        when x"249C" => data_out<= x"8D";
        when x"249D" => data_out<= x"48";
        when x"249E" => data_out<= x"02";
        when x"249F" => data_out<= x"A9";
        when x"24A0" => data_out<= x"01";
        when x"24A1" => data_out<= x"8D";
        when x"24A2" => data_out<= x"47";
        when x"24A3" => data_out<= x"02";
        when x"24A4" => data_out<= x"A2";
        when x"24A5" => data_out<= x"00";
        when x"24A6" => data_out<= x"8A";
        when x"24A7" => data_out<= x"4C";
        when x"24A8" => data_out<= x"2C";
        when x"24A9" => data_out<= x"AF";
        when x"24AA" => data_out<= x"A0";
        when x"24AB" => data_out<= x"02";
        when x"24AC" => data_out<= x"AA";
        when x"24AD" => data_out<= x"B1";
        when x"24AE" => data_out<= x"0C";
        when x"24AF" => data_out<= x"18";
        when x"24B0" => data_out<= x"69";
        when x"24B1" => data_out<= x"01";
        when x"24B2" => data_out<= x"91";
        when x"24B3" => data_out<= x"0C";
        when x"24B4" => data_out<= x"4C";
        when x"24B5" => data_out<= x"F0";
        when x"24B6" => data_out<= x"A3";
        when x"24B7" => data_out<= x"A9";
        when x"24B8" => data_out<= x"03";
        when x"24B9" => data_out<= x"4C";
        when x"24BA" => data_out<= x"2C";
        when x"24BB" => data_out<= x"AF";
        when x"24BC" => data_out<= x"20";
        when x"24BD" => data_out<= x"7B";
        when x"24BE" => data_out<= x"B0";
        when x"24BF" => data_out<= x"20";
        when x"24C0" => data_out<= x"6A";
        when x"24C1" => data_out<= x"AE";
        when x"24C2" => data_out<= x"A9";
        when x"24C3" => data_out<= x"FF";
        when x"24C4" => data_out<= x"20";
        when x"24C5" => data_out<= x"65";
        when x"24C6" => data_out<= x"B0";
        when x"24C7" => data_out<= x"20";
        when x"24C8" => data_out<= x"9A";
        when x"24C9" => data_out<= x"AE";
        when x"24CA" => data_out<= x"20";
        when x"24CB" => data_out<= x"B9";
        when x"24CC" => data_out<= x"A9";
        when x"24CD" => data_out<= x"A9";
        when x"24CE" => data_out<= x"00";
        when x"24CF" => data_out<= x"A0";
        when x"24D0" => data_out<= x"07";
        when x"24D1" => data_out<= x"91";
        when x"24D2" => data_out<= x"0C";
        when x"24D3" => data_out<= x"C9";
        when x"24D4" => data_out<= x"10";
        when x"24D5" => data_out<= x"B0";
        when x"24D6" => data_out<= x"54";
        when x"24D7" => data_out<= x"A2";
        when x"24D8" => data_out<= x"00";
        when x"24D9" => data_out<= x"B1";
        when x"24DA" => data_out<= x"0C";
        when x"24DB" => data_out<= x"20";
        when x"24DC" => data_out<= x"29";
        when x"24DD" => data_out<= x"AE";
        when x"24DE" => data_out<= x"20";
        when x"24DF" => data_out<= x"21";
        when x"24E0" => data_out<= x"AE";
        when x"24E1" => data_out<= x"18";
        when x"24E2" => data_out<= x"69";
        when x"24E3" => data_out<= x"64";
        when x"24E4" => data_out<= x"A8";
        when x"24E5" => data_out<= x"8A";
        when x"24E6" => data_out<= x"69";
        when x"24E7" => data_out<= x"02";
        when x"24E8" => data_out<= x"AA";
        when x"24E9" => data_out<= x"98";
        when x"24EA" => data_out<= x"A0";
        when x"24EB" => data_out<= x"04";
        when x"24EC" => data_out<= x"20";
        when x"24ED" => data_out<= x"C5";
        when x"24EE" => data_out<= x"B0";
        when x"24EF" => data_out<= x"85";
        when x"24F0" => data_out<= x"14";
        when x"24F1" => data_out<= x"86";
        when x"24F2" => data_out<= x"15";
        when x"24F3" => data_out<= x"A0";
        when x"24F4" => data_out<= x"00";
        when x"24F5" => data_out<= x"B1";
        when x"24F6" => data_out<= x"14";
        when x"24F7" => data_out<= x"D0";
        when x"24F8" => data_out<= x"11";
        when x"24F9" => data_out<= x"A0";
        when x"24FA" => data_out<= x"06";
        when x"24FB" => data_out<= x"B1";
        when x"24FC" => data_out<= x"0C";
        when x"24FD" => data_out<= x"C9";
        when x"24FE" => data_out<= x"FF";
        when x"24FF" => data_out<= x"D0";
        when x"2500" => data_out<= x"20";
        when x"2501" => data_out<= x"C8";
        when x"2502" => data_out<= x"B1";
        when x"2503" => data_out<= x"0C";
        when x"2504" => data_out<= x"88";
        when x"2505" => data_out<= x"91";
        when x"2506" => data_out<= x"0C";
        when x"2507" => data_out<= x"4C";
        when x"2508" => data_out<= x"21";
        when x"2509" => data_out<= x"A5";
        when x"250A" => data_out<= x"A0";
        when x"250B" => data_out<= x"07";
        when x"250C" => data_out<= x"20";
        when x"250D" => data_out<= x"93";
        when x"250E" => data_out<= x"B0";
        when x"250F" => data_out<= x"A0";
        when x"2510" => data_out<= x"0D";
        when x"2511" => data_out<= x"20";
        when x"2512" => data_out<= x"4F";
        when x"2513" => data_out<= x"AF";
        when x"2514" => data_out<= x"20";
        when x"2515" => data_out<= x"43";
        when x"2516" => data_out<= x"AB";
        when x"2517" => data_out<= x"AA";
        when x"2518" => data_out<= x"F0";
        when x"2519" => data_out<= x"07";
        when x"251A" => data_out<= x"A2";
        when x"251B" => data_out<= x"00";
        when x"251C" => data_out<= x"A9";
        when x"251D" => data_out<= x"05";
        when x"251E" => data_out<= x"4C";
        when x"251F" => data_out<= x"8D";
        when x"2520" => data_out<= x"A6";
        when x"2521" => data_out<= x"A0";
        when x"2522" => data_out<= x"07";
        when x"2523" => data_out<= x"B1";
        when x"2524" => data_out<= x"0C";
        when x"2525" => data_out<= x"18";
        when x"2526" => data_out<= x"69";
        when x"2527" => data_out<= x"01";
        when x"2528" => data_out<= x"4C";
        when x"2529" => data_out<= x"D1";
        when x"252A" => data_out<= x"A4";
        when x"252B" => data_out<= x"88";
        when x"252C" => data_out<= x"A2";
        when x"252D" => data_out<= x"00";
        when x"252E" => data_out<= x"B1";
        when x"252F" => data_out<= x"0C";
        when x"2530" => data_out<= x"C9";
        when x"2531" => data_out<= x"FF";
        when x"2532" => data_out<= x"D0";
        when x"2533" => data_out<= x"05";
        when x"2534" => data_out<= x"A9";
        when x"2535" => data_out<= x"04";
        when x"2536" => data_out<= x"4C";
        when x"2537" => data_out<= x"8D";
        when x"2538" => data_out<= x"A6";
        when x"2539" => data_out<= x"86";
        when x"253A" => data_out<= x"15";
        when x"253B" => data_out<= x"AD";
        when x"253C" => data_out<= x"5A";
        when x"253D" => data_out<= x"02";
        when x"253E" => data_out<= x"48";
        when x"253F" => data_out<= x"AD";
        when x"2540" => data_out<= x"5B";
        when x"2541" => data_out<= x"02";
        when x"2542" => data_out<= x"05";
        when x"2543" => data_out<= x"15";
        when x"2544" => data_out<= x"AA";
        when x"2545" => data_out<= x"68";
        when x"2546" => data_out<= x"A0";
        when x"2547" => data_out<= x"02";
        when x"2548" => data_out<= x"20";
        when x"2549" => data_out<= x"C5";
        when x"254A" => data_out<= x"B0";
        when x"254B" => data_out<= x"A9";
        when x"254C" => data_out<= x"FF";
        when x"254D" => data_out<= x"18";
        when x"254E" => data_out<= x"A0";
        when x"254F" => data_out<= x"08";
        when x"2550" => data_out<= x"71";
        when x"2551" => data_out<= x"0C";
        when x"2552" => data_out<= x"A9";
        when x"2553" => data_out<= x"01";
        when x"2554" => data_out<= x"C8";
        when x"2555" => data_out<= x"71";
        when x"2556" => data_out<= x"0C";
        when x"2557" => data_out<= x"A2";
        when x"2558" => data_out<= x"00";
        when x"2559" => data_out<= x"4A";
        when x"255A" => data_out<= x"20";
        when x"255B" => data_out<= x"C3";
        when x"255C" => data_out<= x"B0";
        when x"255D" => data_out<= x"C9";
        when x"255E" => data_out<= x"00";
        when x"255F" => data_out<= x"D0";
        when x"2560" => data_out<= x"05";
        when x"2561" => data_out<= x"A9";
        when x"2562" => data_out<= x"01";
        when x"2563" => data_out<= x"20";
        when x"2564" => data_out<= x"C3";
        when x"2565" => data_out<= x"B0";
        when x"2566" => data_out<= x"A0";
        when x"2567" => data_out<= x"06";
        when x"2568" => data_out<= x"B1";
        when x"2569" => data_out<= x"0C";
        when x"256A" => data_out<= x"20";
        when x"256B" => data_out<= x"29";
        when x"256C" => data_out<= x"AE";
        when x"256D" => data_out<= x"20";
        when x"256E" => data_out<= x"21";
        when x"256F" => data_out<= x"AE";
        when x"2570" => data_out<= x"18";
        when x"2571" => data_out<= x"69";
        when x"2572" => data_out<= x"64";
        when x"2573" => data_out<= x"A8";
        when x"2574" => data_out<= x"8A";
        when x"2575" => data_out<= x"69";
        when x"2576" => data_out<= x"02";
        when x"2577" => data_out<= x"AA";
        when x"2578" => data_out<= x"98";
        when x"2579" => data_out<= x"A0";
        when x"257A" => data_out<= x"04";
        when x"257B" => data_out<= x"20";
        when x"257C" => data_out<= x"C5";
        when x"257D" => data_out<= x"B0";
        when x"257E" => data_out<= x"20";
        when x"257F" => data_out<= x"7B";
        when x"2580" => data_out<= x"B0";
        when x"2581" => data_out<= x"A0";
        when x"2582" => data_out<= x"0F";
        when x"2583" => data_out<= x"20";
        when x"2584" => data_out<= x"93";
        when x"2585" => data_out<= x"B0";
        when x"2586" => data_out<= x"A9";
        when x"2587" => data_out<= x"0B";
        when x"2588" => data_out<= x"20";
        when x"2589" => data_out<= x"67";
        when x"258A" => data_out<= x"AB";
        when x"258B" => data_out<= x"A0";
        when x"258C" => data_out<= x"05";
        when x"258D" => data_out<= x"20";
        when x"258E" => data_out<= x"4F";
        when x"258F" => data_out<= x"AF";
        when x"2590" => data_out<= x"85";
        when x"2591" => data_out<= x"14";
        when x"2592" => data_out<= x"86";
        when x"2593" => data_out<= x"15";
        when x"2594" => data_out<= x"A0";
        when x"2595" => data_out<= x"02";
        when x"2596" => data_out<= x"B1";
        when x"2597" => data_out<= x"0C";
        when x"2598" => data_out<= x"A0";
        when x"2599" => data_out<= x"0C";
        when x"259A" => data_out<= x"91";
        when x"259B" => data_out<= x"14";
        when x"259C" => data_out<= x"A0";
        when x"259D" => data_out<= x"05";
        when x"259E" => data_out<= x"20";
        when x"259F" => data_out<= x"4F";
        when x"25A0" => data_out<= x"AF";
        when x"25A1" => data_out<= x"85";
        when x"25A2" => data_out<= x"14";
        when x"25A3" => data_out<= x"86";
        when x"25A4" => data_out<= x"15";
        when x"25A5" => data_out<= x"A0";
        when x"25A6" => data_out<= x"03";
        when x"25A7" => data_out<= x"B1";
        when x"25A8" => data_out<= x"0C";
        when x"25A9" => data_out<= x"A0";
        when x"25AA" => data_out<= x"0D";
        when x"25AB" => data_out<= x"91";
        when x"25AC" => data_out<= x"14";
        when x"25AD" => data_out<= x"A0";
        when x"25AE" => data_out<= x"05";
        when x"25AF" => data_out<= x"20";
        when x"25B0" => data_out<= x"4F";
        when x"25B1" => data_out<= x"AF";
        when x"25B2" => data_out<= x"85";
        when x"25B3" => data_out<= x"14";
        when x"25B4" => data_out<= x"86";
        when x"25B5" => data_out<= x"15";
        when x"25B6" => data_out<= x"A0";
        when x"25B7" => data_out<= x"08";
        when x"25B8" => data_out<= x"B1";
        when x"25B9" => data_out<= x"0C";
        when x"25BA" => data_out<= x"A0";
        when x"25BB" => data_out<= x"0E";
        when x"25BC" => data_out<= x"91";
        when x"25BD" => data_out<= x"14";
        when x"25BE" => data_out<= x"A0";
        when x"25BF" => data_out<= x"05";
        when x"25C0" => data_out<= x"20";
        when x"25C1" => data_out<= x"4F";
        when x"25C2" => data_out<= x"AF";
        when x"25C3" => data_out<= x"85";
        when x"25C4" => data_out<= x"14";
        when x"25C5" => data_out<= x"86";
        when x"25C6" => data_out<= x"15";
        when x"25C7" => data_out<= x"A0";
        when x"25C8" => data_out<= x"09";
        when x"25C9" => data_out<= x"B1";
        when x"25CA" => data_out<= x"0C";
        when x"25CB" => data_out<= x"A0";
        when x"25CC" => data_out<= x"0F";
        when x"25CD" => data_out<= x"91";
        when x"25CE" => data_out<= x"14";
        when x"25CF" => data_out<= x"A0";
        when x"25D0" => data_out<= x"05";
        when x"25D1" => data_out<= x"20";
        when x"25D2" => data_out<= x"4F";
        when x"25D3" => data_out<= x"AF";
        when x"25D4" => data_out<= x"85";
        when x"25D5" => data_out<= x"14";
        when x"25D6" => data_out<= x"86";
        when x"25D7" => data_out<= x"15";
        when x"25D8" => data_out<= x"A0";
        when x"25D9" => data_out<= x"00";
        when x"25DA" => data_out<= x"B1";
        when x"25DB" => data_out<= x"0C";
        when x"25DC" => data_out<= x"A0";
        when x"25DD" => data_out<= x"10";
        when x"25DE" => data_out<= x"91";
        when x"25DF" => data_out<= x"14";
        when x"25E0" => data_out<= x"A0";
        when x"25E1" => data_out<= x"05";
        when x"25E2" => data_out<= x"20";
        when x"25E3" => data_out<= x"4F";
        when x"25E4" => data_out<= x"AF";
        when x"25E5" => data_out<= x"85";
        when x"25E6" => data_out<= x"14";
        when x"25E7" => data_out<= x"86";
        when x"25E8" => data_out<= x"15";
        when x"25E9" => data_out<= x"A0";
        when x"25EA" => data_out<= x"01";
        when x"25EB" => data_out<= x"B1";
        when x"25EC" => data_out<= x"0C";
        when x"25ED" => data_out<= x"A0";
        when x"25EE" => data_out<= x"11";
        when x"25EF" => data_out<= x"91";
        when x"25F0" => data_out<= x"14";
        when x"25F1" => data_out<= x"20";
        when x"25F2" => data_out<= x"4D";
        when x"25F3" => data_out<= x"AF";
        when x"25F4" => data_out<= x"A0";
        when x"25F5" => data_out<= x"02";
        when x"25F6" => data_out<= x"20";
        when x"25F7" => data_out<= x"04";
        when x"25F8" => data_out<= x"AE";
        when x"25F9" => data_out<= x"A0";
        when x"25FA" => data_out<= x"02";
        when x"25FB" => data_out<= x"B1";
        when x"25FC" => data_out<= x"0C";
        when x"25FD" => data_out<= x"8D";
        when x"25FE" => data_out<= x"5A";
        when x"25FF" => data_out<= x"02";
        when x"2600" => data_out<= x"C8";
        when x"2601" => data_out<= x"B1";
        when x"2602" => data_out<= x"0C";
        when x"2603" => data_out<= x"8D";
        when x"2604" => data_out<= x"5B";
        when x"2605" => data_out<= x"02";
        when x"2606" => data_out<= x"20";
        when x"2607" => data_out<= x"37";
        when x"2608" => data_out<= x"AB";
        when x"2609" => data_out<= x"AA";
        when x"260A" => data_out<= x"F0";
        when x"260B" => data_out<= x"07";
        when x"260C" => data_out<= x"A2";
        when x"260D" => data_out<= x"00";
        when x"260E" => data_out<= x"A9";
        when x"260F" => data_out<= x"01";
        when x"2610" => data_out<= x"4C";
        when x"2611" => data_out<= x"8D";
        when x"2612" => data_out<= x"A6";
        when x"2613" => data_out<= x"A9";
        when x"2614" => data_out<= x"54";
        when x"2615" => data_out<= x"A2";
        when x"2616" => data_out<= x"04";
        when x"2617" => data_out<= x"20";
        when x"2618" => data_out<= x"7B";
        when x"2619" => data_out<= x"B0";
        when x"261A" => data_out<= x"A2";
        when x"261B" => data_out<= x"02";
        when x"261C" => data_out<= x"A9";
        when x"261D" => data_out<= x"00";
        when x"261E" => data_out<= x"20";
        when x"261F" => data_out<= x"D2";
        when x"2620" => data_out<= x"AF";
        when x"2621" => data_out<= x"A9";
        when x"2622" => data_out<= x"00";
        when x"2623" => data_out<= x"A0";
        when x"2624" => data_out<= x"07";
        when x"2625" => data_out<= x"91";
        when x"2626" => data_out<= x"0C";
        when x"2627" => data_out<= x"AA";
        when x"2628" => data_out<= x"B1";
        when x"2629" => data_out<= x"0C";
        when x"262A" => data_out<= x"A0";
        when x"262B" => data_out<= x"00";
        when x"262C" => data_out<= x"D1";
        when x"262D" => data_out<= x"0C";
        when x"262E" => data_out<= x"8A";
        when x"262F" => data_out<= x"C8";
        when x"2630" => data_out<= x"F1";
        when x"2631" => data_out<= x"0C";
        when x"2632" => data_out<= x"B0";
        when x"2633" => data_out<= x"51";
        when x"2634" => data_out<= x"A0";
        when x"2635" => data_out<= x"05";
        when x"2636" => data_out<= x"20";
        when x"2637" => data_out<= x"4F";
        when x"2638" => data_out<= x"AF";
        when x"2639" => data_out<= x"85";
        when x"263A" => data_out<= x"14";
        when x"263B" => data_out<= x"86";
        when x"263C" => data_out<= x"15";
        when x"263D" => data_out<= x"A0";
        when x"263E" => data_out<= x"0C";
        when x"263F" => data_out<= x"B1";
        when x"2640" => data_out<= x"14";
        when x"2641" => data_out<= x"20";
        when x"2642" => data_out<= x"79";
        when x"2643" => data_out<= x"B0";
        when x"2644" => data_out<= x"A0";
        when x"2645" => data_out<= x"07";
        when x"2646" => data_out<= x"20";
        when x"2647" => data_out<= x"4F";
        when x"2648" => data_out<= x"AF";
        when x"2649" => data_out<= x"85";
        when x"264A" => data_out<= x"14";
        when x"264B" => data_out<= x"86";
        when x"264C" => data_out<= x"15";
        when x"264D" => data_out<= x"A0";
        when x"264E" => data_out<= x"0D";
        when x"264F" => data_out<= x"B1";
        when x"2650" => data_out<= x"14";
        when x"2651" => data_out<= x"AA";
        when x"2652" => data_out<= x"A9";
        when x"2653" => data_out<= x"00";
        when x"2654" => data_out<= x"20";
        when x"2655" => data_out<= x"43";
        when x"2656" => data_out<= x"B0";
        when x"2657" => data_out<= x"20";
        when x"2658" => data_out<= x"7B";
        when x"2659" => data_out<= x"B0";
        when x"265A" => data_out<= x"A0";
        when x"265B" => data_out<= x"09";
        when x"265C" => data_out<= x"B1";
        when x"265D" => data_out<= x"0C";
        when x"265E" => data_out<= x"20";
        when x"265F" => data_out<= x"E6";
        when x"2660" => data_out<= x"AD";
        when x"2661" => data_out<= x"20";
        when x"2662" => data_out<= x"7B";
        when x"2663" => data_out<= x"B0";
        when x"2664" => data_out<= x"20";
        when x"2665" => data_out<= x"4D";
        when x"2666" => data_out<= x"AF";
        when x"2667" => data_out<= x"20";
        when x"2668" => data_out<= x"4C";
        when x"2669" => data_out<= x"AE";
        when x"266A" => data_out<= x"20";
        when x"266B" => data_out<= x"7E";
        when x"266C" => data_out<= x"AF";
        when x"266D" => data_out<= x"A9";
        when x"266E" => data_out<= x"54";
        when x"266F" => data_out<= x"A2";
        when x"2670" => data_out<= x"04";
        when x"2671" => data_out<= x"20";
        when x"2672" => data_out<= x"B5";
        when x"2673" => data_out<= x"A1";
        when x"2674" => data_out<= x"20";
        when x"2675" => data_out<= x"14";
        when x"2676" => data_out<= x"AF";
        when x"2677" => data_out<= x"A0";
        when x"2678" => data_out<= x"07";
        when x"2679" => data_out<= x"A2";
        when x"267A" => data_out<= x"00";
        when x"267B" => data_out<= x"B1";
        when x"267C" => data_out<= x"0C";
        when x"267D" => data_out<= x"18";
        when x"267E" => data_out<= x"69";
        when x"267F" => data_out<= x"01";
        when x"2680" => data_out<= x"91";
        when x"2681" => data_out<= x"0C";
        when x"2682" => data_out<= x"4C";
        when x"2683" => data_out<= x"28";
        when x"2684" => data_out<= x"A6";
        when x"2685" => data_out<= x"A0";
        when x"2686" => data_out<= x"0B";
        when x"2687" => data_out<= x"20";
        when x"2688" => data_out<= x"4F";
        when x"2689" => data_out<= x"AF";
        when x"268A" => data_out<= x"20";
        when x"268B" => data_out<= x"E0";
        when x"268C" => data_out<= x"A3";
        when x"268D" => data_out<= x"A0";
        when x"268E" => data_out<= x"0C";
        when x"268F" => data_out<= x"4C";
        when x"2690" => data_out<= x"14";
        when x"2691" => data_out<= x"AE";
        when x"2692" => data_out<= x"20";
        when x"2693" => data_out<= x"7B";
        when x"2694" => data_out<= x"B0";
        when x"2695" => data_out<= x"A0";
        when x"2696" => data_out<= x"05";
        when x"2697" => data_out<= x"20";
        when x"2698" => data_out<= x"93";
        when x"2699" => data_out<= x"B0";
        when x"269A" => data_out<= x"20";
        when x"269B" => data_out<= x"77";
        when x"269C" => data_out<= x"B0";
        when x"269D" => data_out<= x"20";
        when x"269E" => data_out<= x"9A";
        when x"269F" => data_out<= x"AE";
        when x"26A0" => data_out<= x"AD";
        when x"26A1" => data_out<= x"47";
        when x"26A2" => data_out<= x"02";
        when x"26A3" => data_out<= x"F0";
        when x"26A4" => data_out<= x"03";
        when x"26A5" => data_out<= x"4C";
        when x"26A6" => data_out<= x"11";
        when x"26A7" => data_out<= x"A8";
        when x"26A8" => data_out<= x"4C";
        when x"26A9" => data_out<= x"36";
        when x"26AA" => data_out<= x"A8";
        when x"26AB" => data_out<= x"AD";
        when x"26AC" => data_out<= x"4A";
        when x"26AD" => data_out<= x"02";
        when x"26AE" => data_out<= x"AE";
        when x"26AF" => data_out<= x"4B";
        when x"26B0" => data_out<= x"02";
        when x"26B1" => data_out<= x"20";
        when x"26B2" => data_out<= x"7B";
        when x"26B3" => data_out<= x"B0";
        when x"26B4" => data_out<= x"AD";
        when x"26B5" => data_out<= x"4F";
        when x"26B6" => data_out<= x"02";
        when x"26B7" => data_out<= x"4A";
        when x"26B8" => data_out<= x"20";
        when x"26B9" => data_out<= x"E6";
        when x"26BA" => data_out<= x"AD";
        when x"26BB" => data_out<= x"A0";
        when x"26BC" => data_out<= x"02";
        when x"26BD" => data_out<= x"20";
        when x"26BE" => data_out<= x"C5";
        when x"26BF" => data_out<= x"B0";
        when x"26C0" => data_out<= x"AD";
        when x"26C1" => data_out<= x"52";
        when x"26C2" => data_out<= x"02";
        when x"26C3" => data_out<= x"C9";
        when x"26C4" => data_out<= x"00";
        when x"26C5" => data_out<= x"AD";
        when x"26C6" => data_out<= x"53";
        when x"26C7" => data_out<= x"02";
        when x"26C8" => data_out<= x"E9";
        when x"26C9" => data_out<= x"02";
        when x"26CA" => data_out<= x"B0";
        when x"26CB" => data_out<= x"13";
        when x"26CC" => data_out<= x"AD";
        when x"26CD" => data_out<= x"50";
        when x"26CE" => data_out<= x"02";
        when x"26CF" => data_out<= x"AE";
        when x"26D0" => data_out<= x"51";
        when x"26D1" => data_out<= x"02";
        when x"26D2" => data_out<= x"20";
        when x"26D3" => data_out<= x"7B";
        when x"26D4" => data_out<= x"B0";
        when x"26D5" => data_out<= x"A0";
        when x"26D6" => data_out<= x"05";
        when x"26D7" => data_out<= x"20";
        when x"26D8" => data_out<= x"4F";
        when x"26D9" => data_out<= x"AF";
        when x"26DA" => data_out<= x"20";
        when x"26DB" => data_out<= x"B6";
        when x"26DC" => data_out<= x"AE";
        when x"26DD" => data_out<= x"F0";
        when x"26DE" => data_out<= x"43";
        when x"26DF" => data_out<= x"AD";
        when x"26E0" => data_out<= x"48";
        when x"26E1" => data_out<= x"02";
        when x"26E2" => data_out<= x"F0";
        when x"26E3" => data_out<= x"18";
        when x"26E4" => data_out<= x"AD";
        when x"26E5" => data_out<= x"50";
        when x"26E6" => data_out<= x"02";
        when x"26E7" => data_out<= x"AE";
        when x"26E8" => data_out<= x"51";
        when x"26E9" => data_out<= x"02";
        when x"26EA" => data_out<= x"20";
        when x"26EB" => data_out<= x"4C";
        when x"26EC" => data_out<= x"AE";
        when x"26ED" => data_out<= x"20";
        when x"26EE" => data_out<= x"7E";
        when x"26EF" => data_out<= x"AF";
        when x"26F0" => data_out<= x"A9";
        when x"26F1" => data_out<= x"54";
        when x"26F2" => data_out<= x"A2";
        when x"26F3" => data_out<= x"04";
        when x"26F4" => data_out<= x"20";
        when x"26F5" => data_out<= x"B5";
        when x"26F6" => data_out<= x"A1";
        when x"26F7" => data_out<= x"A9";
        when x"26F8" => data_out<= x"00";
        when x"26F9" => data_out<= x"8D";
        when x"26FA" => data_out<= x"48";
        when x"26FB" => data_out<= x"02";
        when x"26FC" => data_out<= x"A0";
        when x"26FD" => data_out<= x"03";
        when x"26FE" => data_out<= x"20";
        when x"26FF" => data_out<= x"4F";
        when x"2700" => data_out<= x"AF";
        when x"2701" => data_out<= x"8D";
        when x"2702" => data_out<= x"50";
        when x"2703" => data_out<= x"02";
        when x"2704" => data_out<= x"8E";
        when x"2705" => data_out<= x"51";
        when x"2706" => data_out<= x"02";
        when x"2707" => data_out<= x"20";
        when x"2708" => data_out<= x"4C";
        when x"2709" => data_out<= x"AE";
        when x"270A" => data_out<= x"20";
        when x"270B" => data_out<= x"7E";
        when x"270C" => data_out<= x"AF";
        when x"270D" => data_out<= x"A9";
        when x"270E" => data_out<= x"54";
        when x"270F" => data_out<= x"A2";
        when x"2710" => data_out<= x"04";
        when x"2711" => data_out<= x"20";
        when x"2712" => data_out<= x"0D";
        when x"2713" => data_out<= x"A1";
        when x"2714" => data_out<= x"AC";
        when x"2715" => data_out<= x"4E";
        when x"2716" => data_out<= x"02";
        when x"2717" => data_out<= x"AD";
        when x"2718" => data_out<= x"4F";
        when x"2719" => data_out<= x"02";
        when x"271A" => data_out<= x"29";
        when x"271B" => data_out<= x"01";
        when x"271C" => data_out<= x"8D";
        when x"271D" => data_out<= x"53";
        when x"271E" => data_out<= x"02";
        when x"271F" => data_out<= x"8C";
        when x"2720" => data_out<= x"52";
        when x"2721" => data_out<= x"02";
        when x"2722" => data_out<= x"A9";
        when x"2723" => data_out<= x"00";
        when x"2724" => data_out<= x"38";
        when x"2725" => data_out<= x"ED";
        when x"2726" => data_out<= x"52";
        when x"2727" => data_out<= x"02";
        when x"2728" => data_out<= x"48";
        when x"2729" => data_out<= x"A9";
        when x"272A" => data_out<= x"02";
        when x"272B" => data_out<= x"ED";
        when x"272C" => data_out<= x"53";
        when x"272D" => data_out<= x"02";
        when x"272E" => data_out<= x"AA";
        when x"272F" => data_out<= x"68";
        when x"2730" => data_out<= x"A0";
        when x"2731" => data_out<= x"04";
        when x"2732" => data_out<= x"20";
        when x"2733" => data_out<= x"C5";
        when x"2734" => data_out<= x"B0";
        when x"2735" => data_out<= x"38";
        when x"2736" => data_out<= x"A0";
        when x"2737" => data_out<= x"0A";
        when x"2738" => data_out<= x"F1";
        when x"2739" => data_out<= x"0C";
        when x"273A" => data_out<= x"85";
        when x"273B" => data_out<= x"1C";
        when x"273C" => data_out<= x"8A";
        when x"273D" => data_out<= x"C8";
        when x"273E" => data_out<= x"F1";
        when x"273F" => data_out<= x"0C";
        when x"2740" => data_out<= x"05";
        when x"2741" => data_out<= x"1C";
        when x"2742" => data_out<= x"90";
        when x"2743" => data_out<= x"0A";
        when x"2744" => data_out<= x"F0";
        when x"2745" => data_out<= x"08";
        when x"2746" => data_out<= x"20";
        when x"2747" => data_out<= x"4F";
        when x"2748" => data_out<= x"AF";
        when x"2749" => data_out<= x"A0";
        when x"274A" => data_out<= x"04";
        when x"274B" => data_out<= x"20";
        when x"274C" => data_out<= x"C5";
        when x"274D" => data_out<= x"B0";
        when x"274E" => data_out<= x"A0";
        when x"274F" => data_out<= x"05";
        when x"2750" => data_out<= x"20";
        when x"2751" => data_out<= x"4F";
        when x"2752" => data_out<= x"AF";
        when x"2753" => data_out<= x"18";
        when x"2754" => data_out<= x"6D";
        when x"2755" => data_out<= x"4E";
        when x"2756" => data_out<= x"02";
        when x"2757" => data_out<= x"48";
        when x"2758" => data_out<= x"8A";
        when x"2759" => data_out<= x"6D";
        when x"275A" => data_out<= x"4F";
        when x"275B" => data_out<= x"02";
        when x"275C" => data_out<= x"AA";
        when x"275D" => data_out<= x"68";
        when x"275E" => data_out<= x"38";
        when x"275F" => data_out<= x"ED";
        when x"2760" => data_out<= x"4C";
        when x"2761" => data_out<= x"02";
        when x"2762" => data_out<= x"85";
        when x"2763" => data_out<= x"1C";
        when x"2764" => data_out<= x"8A";
        when x"2765" => data_out<= x"ED";
        when x"2766" => data_out<= x"4D";
        when x"2767" => data_out<= x"02";
        when x"2768" => data_out<= x"05";
        when x"2769" => data_out<= x"1C";
        when x"276A" => data_out<= x"90";
        when x"276B" => data_out<= x"17";
        when x"276C" => data_out<= x"F0";
        when x"276D" => data_out<= x"15";
        when x"276E" => data_out<= x"AD";
        when x"276F" => data_out<= x"4C";
        when x"2770" => data_out<= x"02";
        when x"2771" => data_out<= x"38";
        when x"2772" => data_out<= x"ED";
        when x"2773" => data_out<= x"4E";
        when x"2774" => data_out<= x"02";
        when x"2775" => data_out<= x"48";
        when x"2776" => data_out<= x"AD";
        when x"2777" => data_out<= x"4D";
        when x"2778" => data_out<= x"02";
        when x"2779" => data_out<= x"ED";
        when x"277A" => data_out<= x"4F";
        when x"277B" => data_out<= x"02";
        when x"277C" => data_out<= x"AA";
        when x"277D" => data_out<= x"68";
        when x"277E" => data_out<= x"A0";
        when x"277F" => data_out<= x"04";
        when x"2780" => data_out<= x"20";
        when x"2781" => data_out<= x"C5";
        when x"2782" => data_out<= x"B0";
        when x"2783" => data_out<= x"A2";
        when x"2784" => data_out<= x"00";
        when x"2785" => data_out<= x"8A";
        when x"2786" => data_out<= x"20";
        when x"2787" => data_out<= x"C3";
        when x"2788" => data_out<= x"B0";
        when x"2789" => data_out<= x"20";
        when x"278A" => data_out<= x"7B";
        when x"278B" => data_out<= x"B0";
        when x"278C" => data_out<= x"A0";
        when x"278D" => data_out<= x"07";
        when x"278E" => data_out<= x"20";
        when x"278F" => data_out<= x"4F";
        when x"2790" => data_out<= x"AF";
        when x"2791" => data_out<= x"20";
        when x"2792" => data_out<= x"B6";
        when x"2793" => data_out<= x"AE";
        when x"2794" => data_out<= x"B0";
        when x"2795" => data_out<= x"37";
        when x"2796" => data_out<= x"20";
        when x"2797" => data_out<= x"4D";
        when x"2798" => data_out<= x"AF";
        when x"2799" => data_out<= x"18";
        when x"279A" => data_out<= x"A0";
        when x"279B" => data_out<= x"08";
        when x"279C" => data_out<= x"71";
        when x"279D" => data_out<= x"0C";
        when x"279E" => data_out<= x"85";
        when x"279F" => data_out<= x"0E";
        when x"27A0" => data_out<= x"8A";
        when x"27A1" => data_out<= x"C8";
        when x"27A2" => data_out<= x"71";
        when x"27A3" => data_out<= x"0C";
        when x"27A4" => data_out<= x"85";
        when x"27A5" => data_out<= x"0F";
        when x"27A6" => data_out<= x"20";
        when x"27A7" => data_out<= x"4D";
        when x"27A8" => data_out<= x"AF";
        when x"27A9" => data_out<= x"18";
        when x"27AA" => data_out<= x"6D";
        when x"27AB" => data_out<= x"52";
        when x"27AC" => data_out<= x"02";
        when x"27AD" => data_out<= x"85";
        when x"27AE" => data_out<= x"14";
        when x"27AF" => data_out<= x"8A";
        when x"27B0" => data_out<= x"6D";
        when x"27B1" => data_out<= x"53";
        when x"27B2" => data_out<= x"02";
        when x"27B3" => data_out<= x"18";
        when x"27B4" => data_out<= x"69";
        when x"27B5" => data_out<= x"04";
        when x"27B6" => data_out<= x"85";
        when x"27B7" => data_out<= x"15";
        when x"27B8" => data_out<= x"A0";
        when x"27B9" => data_out<= x"54";
        when x"27BA" => data_out<= x"B1";
        when x"27BB" => data_out<= x"14";
        when x"27BC" => data_out<= x"A0";
        when x"27BD" => data_out<= x"00";
        when x"27BE" => data_out<= x"91";
        when x"27BF" => data_out<= x"0E";
        when x"27C0" => data_out<= x"20";
        when x"27C1" => data_out<= x"4D";
        when x"27C2" => data_out<= x"AF";
        when x"27C3" => data_out<= x"85";
        when x"27C4" => data_out<= x"10";
        when x"27C5" => data_out<= x"86";
        when x"27C6" => data_out<= x"11";
        when x"27C7" => data_out<= x"20";
        when x"27C8" => data_out<= x"E2";
        when x"27C9" => data_out<= x"AE";
        when x"27CA" => data_out<= x"4C";
        when x"27CB" => data_out<= x"86";
        when x"27CC" => data_out<= x"A7";
        when x"27CD" => data_out<= x"A0";
        when x"27CE" => data_out<= x"05";
        when x"27CF" => data_out<= x"20";
        when x"27D0" => data_out<= x"4F";
        when x"27D1" => data_out<= x"AF";
        when x"27D2" => data_out<= x"A0";
        when x"27D3" => data_out<= x"08";
        when x"27D4" => data_out<= x"20";
        when x"27D5" => data_out<= x"04";
        when x"27D6" => data_out<= x"AE";
        when x"27D7" => data_out<= x"A0";
        when x"27D8" => data_out<= x"05";
        when x"27D9" => data_out<= x"20";
        when x"27DA" => data_out<= x"4F";
        when x"27DB" => data_out<= x"AF";
        when x"27DC" => data_out<= x"18";
        when x"27DD" => data_out<= x"6D";
        when x"27DE" => data_out<= x"52";
        when x"27DF" => data_out<= x"02";
        when x"27E0" => data_out<= x"8D";
        when x"27E1" => data_out<= x"52";
        when x"27E2" => data_out<= x"02";
        when x"27E3" => data_out<= x"8A";
        when x"27E4" => data_out<= x"6D";
        when x"27E5" => data_out<= x"53";
        when x"27E6" => data_out<= x"02";
        when x"27E7" => data_out<= x"8D";
        when x"27E8" => data_out<= x"53";
        when x"27E9" => data_out<= x"02";
        when x"27EA" => data_out<= x"A0";
        when x"27EB" => data_out<= x"05";
        when x"27EC" => data_out<= x"20";
        when x"27ED" => data_out<= x"4F";
        when x"27EE" => data_out<= x"AF";
        when x"27EF" => data_out<= x"18";
        when x"27F0" => data_out<= x"6D";
        when x"27F1" => data_out<= x"4E";
        when x"27F2" => data_out<= x"02";
        when x"27F3" => data_out<= x"8D";
        when x"27F4" => data_out<= x"4E";
        when x"27F5" => data_out<= x"02";
        when x"27F6" => data_out<= x"8A";
        when x"27F7" => data_out<= x"6D";
        when x"27F8" => data_out<= x"4F";
        when x"27F9" => data_out<= x"02";
        when x"27FA" => data_out<= x"8D";
        when x"27FB" => data_out<= x"4F";
        when x"27FC" => data_out<= x"02";
        when x"27FD" => data_out<= x"A0";
        when x"27FE" => data_out<= x"05";
        when x"27FF" => data_out<= x"20";
        when x"2800" => data_out<= x"4F";
        when x"2801" => data_out<= x"AF";
        when x"2802" => data_out<= x"A0";
        when x"2803" => data_out<= x"0A";
        when x"2804" => data_out<= x"20";
        when x"2805" => data_out<= x"00";
        when x"2806" => data_out<= x"B1";
        when x"2807" => data_out<= x"A0";
        when x"2808" => data_out<= x"05";
        when x"2809" => data_out<= x"20";
        when x"280A" => data_out<= x"4F";
        when x"280B" => data_out<= x"AF";
        when x"280C" => data_out<= x"A0";
        when x"280D" => data_out<= x"06";
        when x"280E" => data_out<= x"20";
        when x"280F" => data_out<= x"04";
        when x"2810" => data_out<= x"AE";
        when x"2811" => data_out<= x"A0";
        when x"2812" => data_out<= x"0B";
        when x"2813" => data_out<= x"B1";
        when x"2814" => data_out<= x"0C";
        when x"2815" => data_out<= x"88";
        when x"2816" => data_out<= x"11";
        when x"2817" => data_out<= x"0C";
        when x"2818" => data_out<= x"F0";
        when x"2819" => data_out<= x"17";
        when x"281A" => data_out<= x"AD";
        when x"281B" => data_out<= x"4E";
        when x"281C" => data_out<= x"02";
        when x"281D" => data_out<= x"AE";
        when x"281E" => data_out<= x"4F";
        when x"281F" => data_out<= x"02";
        when x"2820" => data_out<= x"20";
        when x"2821" => data_out<= x"7B";
        when x"2822" => data_out<= x"B0";
        when x"2823" => data_out<= x"AD";
        when x"2824" => data_out<= x"4C";
        when x"2825" => data_out<= x"02";
        when x"2826" => data_out<= x"AE";
        when x"2827" => data_out<= x"4D";
        when x"2828" => data_out<= x"02";
        when x"2829" => data_out<= x"20";
        when x"282A" => data_out<= x"B6";
        when x"282B" => data_out<= x"AE";
        when x"282C" => data_out<= x"B0";
        when x"282D" => data_out<= x"03";
        when x"282E" => data_out<= x"4C";
        when x"282F" => data_out<= x"AB";
        when x"2830" => data_out<= x"A6";
        when x"2831" => data_out<= x"A0";
        when x"2832" => data_out<= x"07";
        when x"2833" => data_out<= x"20";
        when x"2834" => data_out<= x"4F";
        when x"2835" => data_out<= x"AF";
        when x"2836" => data_out<= x"A0";
        when x"2837" => data_out<= x"0E";
        when x"2838" => data_out<= x"4C";
        when x"2839" => data_out<= x"14";
        when x"283A" => data_out<= x"AE";
        when x"283B" => data_out<= x"20";
        when x"283C" => data_out<= x"7B";
        when x"283D" => data_out<= x"B0";
        when x"283E" => data_out<= x"A0";
        when x"283F" => data_out<= x"05";
        when x"2840" => data_out<= x"20";
        when x"2841" => data_out<= x"93";
        when x"2842" => data_out<= x"B0";
        when x"2843" => data_out<= x"20";
        when x"2844" => data_out<= x"77";
        when x"2845" => data_out<= x"B0";
        when x"2846" => data_out<= x"20";
        when x"2847" => data_out<= x"8D";
        when x"2848" => data_out<= x"AE";
        when x"2849" => data_out<= x"AD";
        when x"284A" => data_out<= x"47";
        when x"284B" => data_out<= x"02";
        when x"284C" => data_out<= x"F0";
        when x"284D" => data_out<= x"03";
        when x"284E" => data_out<= x"4C";
        when x"284F" => data_out<= x"8F";
        when x"2850" => data_out<= x"A9";
        when x"2851" => data_out<= x"4C";
        when x"2852" => data_out<= x"B4";
        when x"2853" => data_out<= x"A9";
        when x"2854" => data_out<= x"AD";
        when x"2855" => data_out<= x"4A";
        when x"2856" => data_out<= x"02";
        when x"2857" => data_out<= x"AE";
        when x"2858" => data_out<= x"4B";
        when x"2859" => data_out<= x"02";
        when x"285A" => data_out<= x"20";
        when x"285B" => data_out<= x"7B";
        when x"285C" => data_out<= x"B0";
        when x"285D" => data_out<= x"AD";
        when x"285E" => data_out<= x"4F";
        when x"285F" => data_out<= x"02";
        when x"2860" => data_out<= x"4A";
        when x"2861" => data_out<= x"20";
        when x"2862" => data_out<= x"E6";
        when x"2863" => data_out<= x"AD";
        when x"2864" => data_out<= x"20";
        when x"2865" => data_out<= x"C3";
        when x"2866" => data_out<= x"B0";
        when x"2867" => data_out<= x"AD";
        when x"2868" => data_out<= x"52";
        when x"2869" => data_out<= x"02";
        when x"286A" => data_out<= x"C9";
        when x"286B" => data_out<= x"00";
        when x"286C" => data_out<= x"AD";
        when x"286D" => data_out<= x"53";
        when x"286E" => data_out<= x"02";
        when x"286F" => data_out<= x"E9";
        when x"2870" => data_out<= x"02";
        when x"2871" => data_out<= x"B0";
        when x"2872" => data_out<= x"13";
        when x"2873" => data_out<= x"AD";
        when x"2874" => data_out<= x"50";
        when x"2875" => data_out<= x"02";
        when x"2876" => data_out<= x"AE";
        when x"2877" => data_out<= x"51";
        when x"2878" => data_out<= x"02";
        when x"2879" => data_out<= x"20";
        when x"287A" => data_out<= x"7B";
        when x"287B" => data_out<= x"B0";
        when x"287C" => data_out<= x"A0";
        when x"287D" => data_out<= x"03";
        when x"287E" => data_out<= x"20";
        when x"287F" => data_out<= x"4F";
        when x"2880" => data_out<= x"AF";
        when x"2881" => data_out<= x"20";
        when x"2882" => data_out<= x"B6";
        when x"2883" => data_out<= x"AE";
        when x"2884" => data_out<= x"F0";
        when x"2885" => data_out<= x"41";
        when x"2886" => data_out<= x"AD";
        when x"2887" => data_out<= x"48";
        when x"2888" => data_out<= x"02";
        when x"2889" => data_out<= x"F0";
        when x"288A" => data_out<= x"18";
        when x"288B" => data_out<= x"AD";
        when x"288C" => data_out<= x"50";
        when x"288D" => data_out<= x"02";
        when x"288E" => data_out<= x"AE";
        when x"288F" => data_out<= x"51";
        when x"2890" => data_out<= x"02";
        when x"2891" => data_out<= x"20";
        when x"2892" => data_out<= x"4C";
        when x"2893" => data_out<= x"AE";
        when x"2894" => data_out<= x"20";
        when x"2895" => data_out<= x"7E";
        when x"2896" => data_out<= x"AF";
        when x"2897" => data_out<= x"A9";
        when x"2898" => data_out<= x"54";
        when x"2899" => data_out<= x"A2";
        when x"289A" => data_out<= x"04";
        when x"289B" => data_out<= x"20";
        when x"289C" => data_out<= x"B5";
        when x"289D" => data_out<= x"A1";
        when x"289E" => data_out<= x"A9";
        when x"289F" => data_out<= x"00";
        when x"28A0" => data_out<= x"8D";
        when x"28A1" => data_out<= x"48";
        when x"28A2" => data_out<= x"02";
        when x"28A3" => data_out<= x"20";
        when x"28A4" => data_out<= x"4D";
        when x"28A5" => data_out<= x"AF";
        when x"28A6" => data_out<= x"8D";
        when x"28A7" => data_out<= x"50";
        when x"28A8" => data_out<= x"02";
        when x"28A9" => data_out<= x"8E";
        when x"28AA" => data_out<= x"51";
        when x"28AB" => data_out<= x"02";
        when x"28AC" => data_out<= x"20";
        when x"28AD" => data_out<= x"4C";
        when x"28AE" => data_out<= x"AE";
        when x"28AF" => data_out<= x"20";
        when x"28B0" => data_out<= x"7E";
        when x"28B1" => data_out<= x"AF";
        when x"28B2" => data_out<= x"A9";
        when x"28B3" => data_out<= x"54";
        when x"28B4" => data_out<= x"A2";
        when x"28B5" => data_out<= x"04";
        when x"28B6" => data_out<= x"20";
        when x"28B7" => data_out<= x"0D";
        when x"28B8" => data_out<= x"A1";
        when x"28B9" => data_out<= x"AC";
        when x"28BA" => data_out<= x"4E";
        when x"28BB" => data_out<= x"02";
        when x"28BC" => data_out<= x"AD";
        when x"28BD" => data_out<= x"4F";
        when x"28BE" => data_out<= x"02";
        when x"28BF" => data_out<= x"29";
        when x"28C0" => data_out<= x"01";
        when x"28C1" => data_out<= x"8D";
        when x"28C2" => data_out<= x"53";
        when x"28C3" => data_out<= x"02";
        when x"28C4" => data_out<= x"8C";
        when x"28C5" => data_out<= x"52";
        when x"28C6" => data_out<= x"02";
        when x"28C7" => data_out<= x"A9";
        when x"28C8" => data_out<= x"00";
        when x"28C9" => data_out<= x"38";
        when x"28CA" => data_out<= x"ED";
        when x"28CB" => data_out<= x"52";
        when x"28CC" => data_out<= x"02";
        when x"28CD" => data_out<= x"48";
        when x"28CE" => data_out<= x"A9";
        when x"28CF" => data_out<= x"02";
        when x"28D0" => data_out<= x"ED";
        when x"28D1" => data_out<= x"53";
        when x"28D2" => data_out<= x"02";
        when x"28D3" => data_out<= x"AA";
        when x"28D4" => data_out<= x"68";
        when x"28D5" => data_out<= x"A0";
        when x"28D6" => data_out<= x"02";
        when x"28D7" => data_out<= x"20";
        when x"28D8" => data_out<= x"C5";
        when x"28D9" => data_out<= x"B0";
        when x"28DA" => data_out<= x"38";
        when x"28DB" => data_out<= x"A0";
        when x"28DC" => data_out<= x"08";
        when x"28DD" => data_out<= x"F1";
        when x"28DE" => data_out<= x"0C";
        when x"28DF" => data_out<= x"85";
        when x"28E0" => data_out<= x"1C";
        when x"28E1" => data_out<= x"8A";
        when x"28E2" => data_out<= x"C8";
        when x"28E3" => data_out<= x"F1";
        when x"28E4" => data_out<= x"0C";
        when x"28E5" => data_out<= x"05";
        when x"28E6" => data_out<= x"1C";
        when x"28E7" => data_out<= x"90";
        when x"28E8" => data_out<= x"0A";
        when x"28E9" => data_out<= x"F0";
        when x"28EA" => data_out<= x"08";
        when x"28EB" => data_out<= x"20";
        when x"28EC" => data_out<= x"4F";
        when x"28ED" => data_out<= x"AF";
        when x"28EE" => data_out<= x"A0";
        when x"28EF" => data_out<= x"02";
        when x"28F0" => data_out<= x"20";
        when x"28F1" => data_out<= x"C5";
        when x"28F2" => data_out<= x"B0";
        when x"28F3" => data_out<= x"A0";
        when x"28F4" => data_out<= x"03";
        when x"28F5" => data_out<= x"20";
        when x"28F6" => data_out<= x"4F";
        when x"28F7" => data_out<= x"AF";
        when x"28F8" => data_out<= x"18";
        when x"28F9" => data_out<= x"6D";
        when x"28FA" => data_out<= x"4E";
        when x"28FB" => data_out<= x"02";
        when x"28FC" => data_out<= x"48";
        when x"28FD" => data_out<= x"8A";
        when x"28FE" => data_out<= x"6D";
        when x"28FF" => data_out<= x"4F";
        when x"2900" => data_out<= x"02";
        when x"2901" => data_out<= x"AA";
        when x"2902" => data_out<= x"68";
        when x"2903" => data_out<= x"38";
        when x"2904" => data_out<= x"ED";
        when x"2905" => data_out<= x"4C";
        when x"2906" => data_out<= x"02";
        when x"2907" => data_out<= x"85";
        when x"2908" => data_out<= x"1C";
        when x"2909" => data_out<= x"8A";
        when x"290A" => data_out<= x"ED";
        when x"290B" => data_out<= x"4D";
        when x"290C" => data_out<= x"02";
        when x"290D" => data_out<= x"05";
        when x"290E" => data_out<= x"1C";
        when x"290F" => data_out<= x"90";
        when x"2910" => data_out<= x"17";
        when x"2911" => data_out<= x"F0";
        when x"2912" => data_out<= x"15";
        when x"2913" => data_out<= x"AD";
        when x"2914" => data_out<= x"4C";
        when x"2915" => data_out<= x"02";
        when x"2916" => data_out<= x"38";
        when x"2917" => data_out<= x"ED";
        when x"2918" => data_out<= x"4E";
        when x"2919" => data_out<= x"02";
        when x"291A" => data_out<= x"48";
        when x"291B" => data_out<= x"AD";
        when x"291C" => data_out<= x"4D";
        when x"291D" => data_out<= x"02";
        when x"291E" => data_out<= x"ED";
        when x"291F" => data_out<= x"4F";
        when x"2920" => data_out<= x"02";
        when x"2921" => data_out<= x"AA";
        when x"2922" => data_out<= x"68";
        when x"2923" => data_out<= x"A0";
        when x"2924" => data_out<= x"02";
        when x"2925" => data_out<= x"20";
        when x"2926" => data_out<= x"C5";
        when x"2927" => data_out<= x"B0";
        when x"2928" => data_out<= x"AD";
        when x"2929" => data_out<= x"52";
        when x"292A" => data_out<= x"02";
        when x"292B" => data_out<= x"18";
        when x"292C" => data_out<= x"69";
        when x"292D" => data_out<= x"54";
        when x"292E" => data_out<= x"A8";
        when x"292F" => data_out<= x"AD";
        when x"2930" => data_out<= x"53";
        when x"2931" => data_out<= x"02";
        when x"2932" => data_out<= x"69";
        when x"2933" => data_out<= x"04";
        when x"2934" => data_out<= x"AA";
        when x"2935" => data_out<= x"98";
        when x"2936" => data_out<= x"20";
        when x"2937" => data_out<= x"7B";
        when x"2938" => data_out<= x"B0";
        when x"2939" => data_out<= x"A0";
        when x"293A" => data_out<= x"0B";
        when x"293B" => data_out<= x"20";
        when x"293C" => data_out<= x"93";
        when x"293D" => data_out<= x"B0";
        when x"293E" => data_out<= x"A0";
        when x"293F" => data_out<= x"07";
        when x"2940" => data_out<= x"20";
        when x"2941" => data_out<= x"4F";
        when x"2942" => data_out<= x"AF";
        when x"2943" => data_out<= x"20";
        when x"2944" => data_out<= x"96";
        when x"2945" => data_out<= x"AF";
        when x"2946" => data_out<= x"A0";
        when x"2947" => data_out<= x"03";
        when x"2948" => data_out<= x"20";
        when x"2949" => data_out<= x"4F";
        when x"294A" => data_out<= x"AF";
        when x"294B" => data_out<= x"A0";
        when x"294C" => data_out<= x"06";
        when x"294D" => data_out<= x"20";
        when x"294E" => data_out<= x"04";
        when x"294F" => data_out<= x"AE";
        when x"2950" => data_out<= x"A0";
        when x"2951" => data_out<= x"03";
        when x"2952" => data_out<= x"20";
        when x"2953" => data_out<= x"4F";
        when x"2954" => data_out<= x"AF";
        when x"2955" => data_out<= x"18";
        when x"2956" => data_out<= x"6D";
        when x"2957" => data_out<= x"52";
        when x"2958" => data_out<= x"02";
        when x"2959" => data_out<= x"8D";
        when x"295A" => data_out<= x"52";
        when x"295B" => data_out<= x"02";
        when x"295C" => data_out<= x"8A";
        when x"295D" => data_out<= x"6D";
        when x"295E" => data_out<= x"53";
        when x"295F" => data_out<= x"02";
        when x"2960" => data_out<= x"8D";
        when x"2961" => data_out<= x"53";
        when x"2962" => data_out<= x"02";
        when x"2963" => data_out<= x"A0";
        when x"2964" => data_out<= x"03";
        when x"2965" => data_out<= x"20";
        when x"2966" => data_out<= x"4F";
        when x"2967" => data_out<= x"AF";
        when x"2968" => data_out<= x"18";
        when x"2969" => data_out<= x"6D";
        when x"296A" => data_out<= x"4E";
        when x"296B" => data_out<= x"02";
        when x"296C" => data_out<= x"8D";
        when x"296D" => data_out<= x"4E";
        when x"296E" => data_out<= x"02";
        when x"296F" => data_out<= x"8A";
        when x"2970" => data_out<= x"6D";
        when x"2971" => data_out<= x"4F";
        when x"2972" => data_out<= x"02";
        when x"2973" => data_out<= x"8D";
        when x"2974" => data_out<= x"4F";
        when x"2975" => data_out<= x"02";
        when x"2976" => data_out<= x"A0";
        when x"2977" => data_out<= x"03";
        when x"2978" => data_out<= x"20";
        when x"2979" => data_out<= x"4F";
        when x"297A" => data_out<= x"AF";
        when x"297B" => data_out<= x"A0";
        when x"297C" => data_out<= x"08";
        when x"297D" => data_out<= x"20";
        when x"297E" => data_out<= x"00";
        when x"297F" => data_out<= x"B1";
        when x"2980" => data_out<= x"A0";
        when x"2981" => data_out<= x"03";
        when x"2982" => data_out<= x"20";
        when x"2983" => data_out<= x"4F";
        when x"2984" => data_out<= x"AF";
        when x"2985" => data_out<= x"A0";
        when x"2986" => data_out<= x"04";
        when x"2987" => data_out<= x"20";
        when x"2988" => data_out<= x"04";
        when x"2989" => data_out<= x"AE";
        when x"298A" => data_out<= x"A9";
        when x"298B" => data_out<= x"01";
        when x"298C" => data_out<= x"8D";
        when x"298D" => data_out<= x"48";
        when x"298E" => data_out<= x"02";
        when x"298F" => data_out<= x"A0";
        when x"2990" => data_out<= x"09";
        when x"2991" => data_out<= x"B1";
        when x"2992" => data_out<= x"0C";
        when x"2993" => data_out<= x"88";
        when x"2994" => data_out<= x"11";
        when x"2995" => data_out<= x"0C";
        when x"2996" => data_out<= x"F0";
        when x"2997" => data_out<= x"17";
        when x"2998" => data_out<= x"AD";
        when x"2999" => data_out<= x"4E";
        when x"299A" => data_out<= x"02";
        when x"299B" => data_out<= x"AE";
        when x"299C" => data_out<= x"4F";
        when x"299D" => data_out<= x"02";
        when x"299E" => data_out<= x"20";
        when x"299F" => data_out<= x"7B";
        when x"29A0" => data_out<= x"B0";
        when x"29A1" => data_out<= x"AD";
        when x"29A2" => data_out<= x"4C";
        when x"29A3" => data_out<= x"02";
        when x"29A4" => data_out<= x"AE";
        when x"29A5" => data_out<= x"4D";
        when x"29A6" => data_out<= x"02";
        when x"29A7" => data_out<= x"20";
        when x"29A8" => data_out<= x"B6";
        when x"29A9" => data_out<= x"AE";
        when x"29AA" => data_out<= x"B0";
        when x"29AB" => data_out<= x"03";
        when x"29AC" => data_out<= x"4C";
        when x"29AD" => data_out<= x"54";
        when x"29AE" => data_out<= x"A8";
        when x"29AF" => data_out<= x"A0";
        when x"29B0" => data_out<= x"05";
        when x"29B1" => data_out<= x"20";
        when x"29B2" => data_out<= x"4F";
        when x"29B3" => data_out<= x"AF";
        when x"29B4" => data_out<= x"A0";
        when x"29B5" => data_out<= x"0C";
        when x"29B6" => data_out<= x"4C";
        when x"29B7" => data_out<= x"14";
        when x"29B8" => data_out<= x"AE";
        when x"29B9" => data_out<= x"AD";
        when x"29BA" => data_out<= x"47";
        when x"29BB" => data_out<= x"02";
        when x"29BC" => data_out<= x"F0";
        when x"29BD" => data_out<= x"20";
        when x"29BE" => data_out<= x"AD";
        when x"29BF" => data_out<= x"48";
        when x"29C0" => data_out<= x"02";
        when x"29C1" => data_out<= x"F0";
        when x"29C2" => data_out<= x"15";
        when x"29C3" => data_out<= x"AD";
        when x"29C4" => data_out<= x"50";
        when x"29C5" => data_out<= x"02";
        when x"29C6" => data_out<= x"AE";
        when x"29C7" => data_out<= x"51";
        when x"29C8" => data_out<= x"02";
        when x"29C9" => data_out<= x"20";
        when x"29CA" => data_out<= x"4C";
        when x"29CB" => data_out<= x"AE";
        when x"29CC" => data_out<= x"20";
        when x"29CD" => data_out<= x"7E";
        when x"29CE" => data_out<= x"AF";
        when x"29CF" => data_out<= x"A9";
        when x"29D0" => data_out<= x"54";
        when x"29D1" => data_out<= x"A2";
        when x"29D2" => data_out<= x"04";
        when x"29D3" => data_out<= x"20";
        when x"29D4" => data_out<= x"B5";
        when x"29D5" => data_out<= x"A1";
        when x"29D6" => data_out<= x"A9";
        when x"29D7" => data_out<= x"00";
        when x"29D8" => data_out<= x"8D";
        when x"29D9" => data_out<= x"47";
        when x"29DA" => data_out<= x"02";
        when x"29DB" => data_out<= x"8D";
        when x"29DC" => data_out<= x"48";
        when x"29DD" => data_out<= x"02";
        when x"29DE" => data_out<= x"60";
        when x"29DF" => data_out<= x"20";
        when x"29E0" => data_out<= x"7B";
        when x"29E1" => data_out<= x"B0";
        when x"29E2" => data_out<= x"20";
        when x"29E3" => data_out<= x"80";
        when x"29E4" => data_out<= x"AE";
        when x"29E5" => data_out<= x"20";
        when x"29E6" => data_out<= x"B9";
        when x"29E7" => data_out<= x"A9";
        when x"29E8" => data_out<= x"A9";
        when x"29E9" => data_out<= x"00";
        when x"29EA" => data_out<= x"A0";
        when x"29EB" => data_out<= x"02";
        when x"29EC" => data_out<= x"91";
        when x"29ED" => data_out<= x"0C";
        when x"29EE" => data_out<= x"AA";
        when x"29EF" => data_out<= x"B1";
        when x"29F0" => data_out<= x"0C";
        when x"29F1" => data_out<= x"C9";
        when x"29F2" => data_out<= x"10";
        when x"29F3" => data_out<= x"B0";
        when x"29F4" => data_out<= x"57";
        when x"29F5" => data_out<= x"20";
        when x"29F6" => data_out<= x"29";
        when x"29F7" => data_out<= x"AE";
        when x"29F8" => data_out<= x"20";
        when x"29F9" => data_out<= x"21";
        when x"29FA" => data_out<= x"AE";
        when x"29FB" => data_out<= x"18";
        when x"29FC" => data_out<= x"69";
        when x"29FD" => data_out<= x"64";
        when x"29FE" => data_out<= x"A8";
        when x"29FF" => data_out<= x"8A";
        when x"2A00" => data_out<= x"69";
        when x"2A01" => data_out<= x"02";
        when x"2A02" => data_out<= x"AA";
        when x"2A03" => data_out<= x"98";
        when x"2A04" => data_out<= x"20";
        when x"2A05" => data_out<= x"C3";
        when x"2A06" => data_out<= x"B0";
        when x"2A07" => data_out<= x"85";
        when x"2A08" => data_out<= x"14";
        when x"2A09" => data_out<= x"86";
        when x"2A0A" => data_out<= x"15";
        when x"2A0B" => data_out<= x"A0";
        when x"2A0C" => data_out<= x"00";
        when x"2A0D" => data_out<= x"B1";
        when x"2A0E" => data_out<= x"14";
        when x"2A0F" => data_out<= x"F0";
        when x"2A10" => data_out<= x"2E";
        when x"2A11" => data_out<= x"20";
        when x"2A12" => data_out<= x"91";
        when x"2A13" => data_out<= x"B0";
        when x"2A14" => data_out<= x"A0";
        when x"2A15" => data_out<= x"06";
        when x"2A16" => data_out<= x"20";
        when x"2A17" => data_out<= x"4F";
        when x"2A18" => data_out<= x"AF";
        when x"2A19" => data_out<= x"20";
        when x"2A1A" => data_out<= x"43";
        when x"2A1B" => data_out<= x"AB";
        when x"2A1C" => data_out<= x"AA";
        when x"2A1D" => data_out<= x"F0";
        when x"2A1E" => data_out<= x"20";
        when x"2A1F" => data_out<= x"20";
        when x"2A20" => data_out<= x"4D";
        when x"2A21" => data_out<= x"AF";
        when x"2A22" => data_out<= x"85";
        when x"2A23" => data_out<= x"14";
        when x"2A24" => data_out<= x"86";
        when x"2A25" => data_out<= x"15";
        when x"2A26" => data_out<= x"A9";
        when x"2A27" => data_out<= x"00";
        when x"2A28" => data_out<= x"A8";
        when x"2A29" => data_out<= x"91";
        when x"2A2A" => data_out<= x"14";
        when x"2A2B" => data_out<= x"20";
        when x"2A2C" => data_out<= x"37";
        when x"2A2D" => data_out<= x"AB";
        when x"2A2E" => data_out<= x"86";
        when x"2A2F" => data_out<= x"1C";
        when x"2A30" => data_out<= x"05";
        when x"2A31" => data_out<= x"1C";
        when x"2A32" => data_out<= x"F0";
        when x"2A33" => data_out<= x"07";
        when x"2A34" => data_out<= x"A2";
        when x"2A35" => data_out<= x"00";
        when x"2A36" => data_out<= x"A9";
        when x"2A37" => data_out<= x"01";
        when x"2A38" => data_out<= x"4C";
        when x"2A39" => data_out<= x"2C";
        when x"2A3A" => data_out<= x"AF";
        when x"2A3B" => data_out<= x"AA";
        when x"2A3C" => data_out<= x"4C";
        when x"2A3D" => data_out<= x"2C";
        when x"2A3E" => data_out<= x"AF";
        when x"2A3F" => data_out<= x"A0";
        when x"2A40" => data_out<= x"02";
        when x"2A41" => data_out<= x"AA";
        when x"2A42" => data_out<= x"B1";
        when x"2A43" => data_out<= x"0C";
        when x"2A44" => data_out<= x"18";
        when x"2A45" => data_out<= x"69";
        when x"2A46" => data_out<= x"01";
        when x"2A47" => data_out<= x"91";
        when x"2A48" => data_out<= x"0C";
        when x"2A49" => data_out<= x"4C";
        when x"2A4A" => data_out<= x"EF";
        when x"2A4B" => data_out<= x"A9";
        when x"2A4C" => data_out<= x"A9";
        when x"2A4D" => data_out<= x"03";
        when x"2A4E" => data_out<= x"4C";
        when x"2A4F" => data_out<= x"2C";
        when x"2A50" => data_out<= x"AF";
        when x"2A51" => data_out<= x"20";
        when x"2A52" => data_out<= x"7B";
        when x"2A53" => data_out<= x"B0";
        when x"2A54" => data_out<= x"20";
        when x"2A55" => data_out<= x"80";
        when x"2A56" => data_out<= x"AE";
        when x"2A57" => data_out<= x"A0";
        when x"2A58" => data_out<= x"05";
        when x"2A59" => data_out<= x"B1";
        when x"2A5A" => data_out<= x"0C";
        when x"2A5B" => data_out<= x"C9";
        when x"2A5C" => data_out<= x"10";
        when x"2A5D" => data_out<= x"A2";
        when x"2A5E" => data_out<= x"00";
        when x"2A5F" => data_out<= x"90";
        when x"2A60" => data_out<= x"05";
        when x"2A61" => data_out<= x"A9";
        when x"2A62" => data_out<= x"03";
        when x"2A63" => data_out<= x"4C";
        when x"2A64" => data_out<= x"31";
        when x"2A65" => data_out<= x"AF";
        when x"2A66" => data_out<= x"B1";
        when x"2A67" => data_out<= x"0C";
        when x"2A68" => data_out<= x"20";
        when x"2A69" => data_out<= x"29";
        when x"2A6A" => data_out<= x"AE";
        when x"2A6B" => data_out<= x"20";
        when x"2A6C" => data_out<= x"21";
        when x"2A6D" => data_out<= x"AE";
        when x"2A6E" => data_out<= x"18";
        when x"2A6F" => data_out<= x"69";
        when x"2A70" => data_out<= x"64";
        when x"2A71" => data_out<= x"A8";
        when x"2A72" => data_out<= x"8A";
        when x"2A73" => data_out<= x"69";
        when x"2A74" => data_out<= x"02";
        when x"2A75" => data_out<= x"AA";
        when x"2A76" => data_out<= x"98";
        when x"2A77" => data_out<= x"A0";
        when x"2A78" => data_out<= x"01";
        when x"2A79" => data_out<= x"20";
        when x"2A7A" => data_out<= x"C5";
        when x"2A7B" => data_out<= x"B0";
        when x"2A7C" => data_out<= x"85";
        when x"2A7D" => data_out<= x"14";
        when x"2A7E" => data_out<= x"86";
        when x"2A7F" => data_out<= x"15";
        when x"2A80" => data_out<= x"A0";
        when x"2A81" => data_out<= x"00";
        when x"2A82" => data_out<= x"B1";
        when x"2A83" => data_out<= x"14";
        when x"2A84" => data_out<= x"D0";
        when x"2A85" => data_out<= x"06";
        when x"2A86" => data_out<= x"AA";
        when x"2A87" => data_out<= x"A9";
        when x"2A88" => data_out<= x"03";
        when x"2A89" => data_out<= x"4C";
        when x"2A8A" => data_out<= x"31";
        when x"2A8B" => data_out<= x"AF";
        when x"2A8C" => data_out<= x"98";
        when x"2A8D" => data_out<= x"91";
        when x"2A8E" => data_out<= x"0C";
        when x"2A8F" => data_out<= x"C9";
        when x"2A90" => data_out<= x"0B";
        when x"2A91" => data_out<= x"B0";
        when x"2A92" => data_out<= x"44";
        when x"2A93" => data_out<= x"A0";
        when x"2A94" => data_out<= x"02";
        when x"2A95" => data_out<= x"20";
        when x"2A96" => data_out<= x"4F";
        when x"2A97" => data_out<= x"AF";
        when x"2A98" => data_out<= x"85";
        when x"2A99" => data_out<= x"14";
        when x"2A9A" => data_out<= x"86";
        when x"2A9B" => data_out<= x"15";
        when x"2A9C" => data_out<= x"A0";
        when x"2A9D" => data_out<= x"00";
        when x"2A9E" => data_out<= x"B1";
        when x"2A9F" => data_out<= x"0C";
        when x"2AA0" => data_out<= x"A8";
        when x"2AA1" => data_out<= x"B1";
        when x"2AA2" => data_out<= x"14";
        when x"2AA3" => data_out<= x"F0";
        when x"2AA4" => data_out<= x"32";
        when x"2AA5" => data_out<= x"A2";
        when x"2AA6" => data_out<= x"00";
        when x"2AA7" => data_out<= x"A1";
        when x"2AA8" => data_out<= x"0C";
        when x"2AA9" => data_out<= x"18";
        when x"2AAA" => data_out<= x"A0";
        when x"2AAB" => data_out<= x"03";
        when x"2AAC" => data_out<= x"71";
        when x"2AAD" => data_out<= x"0C";
        when x"2AAE" => data_out<= x"48";
        when x"2AAF" => data_out<= x"8A";
        when x"2AB0" => data_out<= x"C8";
        when x"2AB1" => data_out<= x"71";
        when x"2AB2" => data_out<= x"0C";
        when x"2AB3" => data_out<= x"AA";
        when x"2AB4" => data_out<= x"68";
        when x"2AB5" => data_out<= x"20";
        when x"2AB6" => data_out<= x"7B";
        when x"2AB7" => data_out<= x"B0";
        when x"2AB8" => data_out<= x"A0";
        when x"2AB9" => data_out<= x"04";
        when x"2ABA" => data_out<= x"20";
        when x"2ABB" => data_out<= x"4F";
        when x"2ABC" => data_out<= x"AF";
        when x"2ABD" => data_out<= x"85";
        when x"2ABE" => data_out<= x"14";
        when x"2ABF" => data_out<= x"86";
        when x"2AC0" => data_out<= x"15";
        when x"2AC1" => data_out<= x"A0";
        when x"2AC2" => data_out<= x"02";
        when x"2AC3" => data_out<= x"B1";
        when x"2AC4" => data_out<= x"0C";
        when x"2AC5" => data_out<= x"A8";
        when x"2AC6" => data_out<= x"B1";
        when x"2AC7" => data_out<= x"14";
        when x"2AC8" => data_out<= x"A0";
        when x"2AC9" => data_out<= x"00";
        when x"2ACA" => data_out<= x"20";
        when x"2ACB" => data_out<= x"AD";
        when x"2ACC" => data_out<= x"B0";
        when x"2ACD" => data_out<= x"A0";
        when x"2ACE" => data_out<= x"00";
        when x"2ACF" => data_out<= x"B1";
        when x"2AD0" => data_out<= x"0C";
        when x"2AD1" => data_out<= x"18";
        when x"2AD2" => data_out<= x"69";
        when x"2AD3" => data_out<= x"01";
        when x"2AD4" => data_out<= x"4C";
        when x"2AD5" => data_out<= x"8D";
        when x"2AD6" => data_out<= x"AA";
        when x"2AD7" => data_out<= x"A2";
        when x"2AD8" => data_out<= x"00";
        when x"2AD9" => data_out<= x"A1";
        when x"2ADA" => data_out<= x"0C";
        when x"2ADB" => data_out<= x"18";
        when x"2ADC" => data_out<= x"A0";
        when x"2ADD" => data_out<= x"03";
        when x"2ADE" => data_out<= x"71";
        when x"2ADF" => data_out<= x"0C";
        when x"2AE0" => data_out<= x"85";
        when x"2AE1" => data_out<= x"14";
        when x"2AE2" => data_out<= x"8A";
        when x"2AE3" => data_out<= x"C8";
        when x"2AE4" => data_out<= x"71";
        when x"2AE5" => data_out<= x"0C";
        when x"2AE6" => data_out<= x"85";
        when x"2AE7" => data_out<= x"15";
        when x"2AE8" => data_out<= x"8A";
        when x"2AE9" => data_out<= x"A8";
        when x"2AEA" => data_out<= x"91";
        when x"2AEB" => data_out<= x"14";
        when x"2AEC" => data_out<= x"A0";
        when x"2AED" => data_out<= x"06";
        when x"2AEE" => data_out<= x"20";
        when x"2AEF" => data_out<= x"93";
        when x"2AF0" => data_out<= x"B0";
        when x"2AF1" => data_out<= x"A0";
        when x"2AF2" => data_out<= x"04";
        when x"2AF3" => data_out<= x"20";
        when x"2AF4" => data_out<= x"4F";
        when x"2AF5" => data_out<= x"AF";
        when x"2AF6" => data_out<= x"85";
        when x"2AF7" => data_out<= x"14";
        when x"2AF8" => data_out<= x"86";
        when x"2AF9" => data_out<= x"15";
        when x"2AFA" => data_out<= x"A0";
        when x"2AFB" => data_out<= x"0E";
        when x"2AFC" => data_out<= x"B1";
        when x"2AFD" => data_out<= x"14";
        when x"2AFE" => data_out<= x"20";
        when x"2AFF" => data_out<= x"79";
        when x"2B00" => data_out<= x"B0";
        when x"2B01" => data_out<= x"A0";
        when x"2B02" => data_out<= x"06";
        when x"2B03" => data_out<= x"20";
        when x"2B04" => data_out<= x"4F";
        when x"2B05" => data_out<= x"AF";
        when x"2B06" => data_out<= x"85";
        when x"2B07" => data_out<= x"14";
        when x"2B08" => data_out<= x"86";
        when x"2B09" => data_out<= x"15";
        when x"2B0A" => data_out<= x"A0";
        when x"2B0B" => data_out<= x"0F";
        when x"2B0C" => data_out<= x"B1";
        when x"2B0D" => data_out<= x"14";
        when x"2B0E" => data_out<= x"AA";
        when x"2B0F" => data_out<= x"A9";
        when x"2B10" => data_out<= x"00";
        when x"2B11" => data_out<= x"20";
        when x"2B12" => data_out<= x"43";
        when x"2B13" => data_out<= x"B0";
        when x"2B14" => data_out<= x"A0";
        when x"2B15" => data_out<= x"0C";
        when x"2B16" => data_out<= x"20";
        when x"2B17" => data_out<= x"CE";
        when x"2B18" => data_out<= x"B0";
        when x"2B19" => data_out<= x"A0";
        when x"2B1A" => data_out<= x"04";
        when x"2B1B" => data_out<= x"20";
        when x"2B1C" => data_out<= x"4F";
        when x"2B1D" => data_out<= x"AF";
        when x"2B1E" => data_out<= x"85";
        when x"2B1F" => data_out<= x"14";
        when x"2B20" => data_out<= x"86";
        when x"2B21" => data_out<= x"15";
        when x"2B22" => data_out<= x"A0";
        when x"2B23" => data_out<= x"05";
        when x"2B24" => data_out<= x"B1";
        when x"2B25" => data_out<= x"0C";
        when x"2B26" => data_out<= x"A0";
        when x"2B27" => data_out<= x"0E";
        when x"2B28" => data_out<= x"91";
        when x"2B29" => data_out<= x"14";
        when x"2B2A" => data_out<= x"A2";
        when x"2B2B" => data_out<= x"00";
        when x"2B2C" => data_out<= x"8A";
        when x"2B2D" => data_out<= x"4C";
        when x"2B2E" => data_out<= x"31";
        when x"2B2F" => data_out<= x"AF";
        when x"2B30" => data_out<= x"AD";
        when x"2B31" => data_out<= x"4C";
        when x"2B32" => data_out<= x"02";
        when x"2B33" => data_out<= x"AE";
        when x"2B34" => data_out<= x"4D";
        when x"2B35" => data_out<= x"02";
        when x"2B36" => data_out<= x"60";
        when x"2B37" => data_out<= x"A2";
        when x"2B38" => data_out<= x"00";
        when x"2B39" => data_out<= x"20";
        when x"2B3A" => data_out<= x"75";
        when x"2B3B" => data_out<= x"AF";
        when x"2B3C" => data_out<= x"A9";
        when x"2B3D" => data_out<= x"54";
        when x"2B3E" => data_out<= x"A2";
        when x"2B3F" => data_out<= x"02";
        when x"2B40" => data_out<= x"4C";
        when x"2B41" => data_out<= x"B5";
        when x"2B42" => data_out<= x"A1";
        when x"2B43" => data_out<= x"85";
        when x"2B44" => data_out<= x"16";
        when x"2B45" => data_out<= x"86";
        when x"2B46" => data_out<= x"17";
        when x"2B47" => data_out<= x"20";
        when x"2B48" => data_out<= x"0C";
        when x"2B49" => data_out<= x"AF";
        when x"2B4A" => data_out<= x"85";
        when x"2B4B" => data_out<= x"14";
        when x"2B4C" => data_out<= x"86";
        when x"2B4D" => data_out<= x"15";
        when x"2B4E" => data_out<= x"A0";
        when x"2B4F" => data_out<= x"00";
        when x"2B50" => data_out<= x"B1";
        when x"2B51" => data_out<= x"14";
        when x"2B52" => data_out<= x"D1";
        when x"2B53" => data_out<= x"16";
        when x"2B54" => data_out<= x"D0";
        when x"2B55" => data_out<= x"07";
        when x"2B56" => data_out<= x"C9";
        when x"2B57" => data_out<= x"00";
        when x"2B58" => data_out<= x"F0";
        when x"2B59" => data_out<= x"08";
        when x"2B5A" => data_out<= x"C8";
        when x"2B5B" => data_out<= x"D0";
        when x"2B5C" => data_out<= x"F3";
        when x"2B5D" => data_out<= x"A9";
        when x"2B5E" => data_out<= x"00";
        when x"2B5F" => data_out<= x"A2";
        when x"2B60" => data_out<= x"00";
        when x"2B61" => data_out<= x"60";
        when x"2B62" => data_out<= x"A9";
        when x"2B63" => data_out<= x"01";
        when x"2B64" => data_out<= x"A2";
        when x"2B65" => data_out<= x"00";
        when x"2B66" => data_out<= x"60";
        when x"2B67" => data_out<= x"85";
        when x"2B68" => data_out<= x"1C";
        when x"2B69" => data_out<= x"20";
        when x"2B6A" => data_out<= x"0C";
        when x"2B6B" => data_out<= x"AF";
        when x"2B6C" => data_out<= x"85";
        when x"2B6D" => data_out<= x"16";
        when x"2B6E" => data_out<= x"86";
        when x"2B6F" => data_out<= x"17";
        when x"2B70" => data_out<= x"20";
        when x"2B71" => data_out<= x"0C";
        when x"2B72" => data_out<= x"AF";
        when x"2B73" => data_out<= x"85";
        when x"2B74" => data_out<= x"14";
        when x"2B75" => data_out<= x"86";
        when x"2B76" => data_out<= x"15";
        when x"2B77" => data_out<= x"A0";
        when x"2B78" => data_out<= x"00";
        when x"2B79" => data_out<= x"A5";
        when x"2B7A" => data_out<= x"1C";
        when x"2B7B" => data_out<= x"F0";
        when x"2B7C" => data_out<= x"0B";
        when x"2B7D" => data_out<= x"C6";
        when x"2B7E" => data_out<= x"1C";
        when x"2B7F" => data_out<= x"B1";
        when x"2B80" => data_out<= x"16";
        when x"2B81" => data_out<= x"F0";
        when x"2B82" => data_out<= x"05";
        when x"2B83" => data_out<= x"91";
        when x"2B84" => data_out<= x"14";
        when x"2B85" => data_out<= x"C8";
        when x"2B86" => data_out<= x"D0";
        when x"2B87" => data_out<= x"F1";
        when x"2B88" => data_out<= x"A9";
        when x"2B89" => data_out<= x"00";
        when x"2B8A" => data_out<= x"91";
        when x"2B8B" => data_out<= x"14";
        when x"2B8C" => data_out<= x"60";
        when x"2B8D" => data_out<= x"A5";
        when x"2B8E" => data_out<= x"0C";
        when x"2B8F" => data_out<= x"48";
        when x"2B90" => data_out<= x"A5";
        when x"2B91" => data_out<= x"0D";
        when x"2B92" => data_out<= x"48";
        when x"2B93" => data_out<= x"A9";
        when x"2B94" => data_out<= x"00";
        when x"2B95" => data_out<= x"85";
        when x"2B96" => data_out<= x"0C";
        when x"2B97" => data_out<= x"A9";
        when x"2B98" => data_out<= x"3F";
        when x"2B99" => data_out<= x"85";
        when x"2B9A" => data_out<= x"0D";
        when x"2B9B" => data_out<= x"38";
        when x"2B9C" => data_out<= x"A5";
        when x"2B9D" => data_out<= x"0C";
        when x"2B9E" => data_out<= x"E9";
        when x"2B9F" => data_out<= x"02";
        when x"2BA0" => data_out<= x"85";
        when x"2BA1" => data_out<= x"0C";
        when x"2BA2" => data_out<= x"B0";
        when x"2BA3" => data_out<= x"02";
        when x"2BA4" => data_out<= x"C6";
        when x"2BA5" => data_out<= x"0D";
        when x"2BA6" => data_out<= x"A0";
        when x"2BA7" => data_out<= x"00";
        when x"2BA8" => data_out<= x"A5";
        when x"2BA9" => data_out<= x"F0";
        when x"2BAA" => data_out<= x"91";
        when x"2BAB" => data_out<= x"0C";
        when x"2BAC" => data_out<= x"C8";
        when x"2BAD" => data_out<= x"A5";
        when x"2BAE" => data_out<= x"F1";
        when x"2BAF" => data_out<= x"91";
        when x"2BB0" => data_out<= x"0C";
        when x"2BB1" => data_out<= x"A5";
        when x"2BB2" => data_out<= x"F2";
        when x"2BB3" => data_out<= x"A6";
        when x"2BB4" => data_out<= x"F3";
        when x"2BB5" => data_out<= x"20";
        when x"2BB6" => data_out<= x"92";
        when x"2BB7" => data_out<= x"A6";
        when x"2BB8" => data_out<= x"85";
        when x"2BB9" => data_out<= x"F2";
        when x"2BBA" => data_out<= x"86";
        when x"2BBB" => data_out<= x"F3";
        when x"2BBC" => data_out<= x"68";
        when x"2BBD" => data_out<= x"85";
        when x"2BBE" => data_out<= x"0D";
        when x"2BBF" => data_out<= x"68";
        when x"2BC0" => data_out<= x"85";
        when x"2BC1" => data_out<= x"0C";
        when x"2BC2" => data_out<= x"A5";
        when x"2BC3" => data_out<= x"F2";
        when x"2BC4" => data_out<= x"A6";
        when x"2BC5" => data_out<= x"F3";
        when x"2BC6" => data_out<= x"60";
        when x"2BC7" => data_out<= x"20";
        when x"2BC8" => data_out<= x"7B";
        when x"2BC9" => data_out<= x"B0";
        when x"2BCA" => data_out<= x"20";
        when x"2BCB" => data_out<= x"91";
        when x"2BCC" => data_out<= x"B0";
        when x"2BCD" => data_out<= x"A9";
        when x"2BCE" => data_out<= x"01";
        when x"2BCF" => data_out<= x"20";
        when x"2BD0" => data_out<= x"65";
        when x"2BD1" => data_out<= x"B0";
        when x"2BD2" => data_out<= x"20";
        when x"2BD3" => data_out<= x"77";
        when x"2BD4" => data_out<= x"B0";
        when x"2BD5" => data_out<= x"A0";
        when x"2BD6" => data_out<= x"09";
        when x"2BD7" => data_out<= x"20";
        when x"2BD8" => data_out<= x"13";
        when x"2BD9" => data_out<= x"B1";
        when x"2BDA" => data_out<= x"A9";
        when x"2BDB" => data_out<= x"00";
        when x"2BDC" => data_out<= x"A0";
        when x"2BDD" => data_out<= x"02";
        when x"2BDE" => data_out<= x"91";
        when x"2BDF" => data_out<= x"0C";
        when x"2BE0" => data_out<= x"C9";
        when x"2BE1" => data_out<= x"3C";
        when x"2BE2" => data_out<= x"B0";
        when x"2BE3" => data_out<= x"60";
        when x"2BE4" => data_out<= x"A9";
        when x"2BE5" => data_out<= x"15";
        when x"2BE6" => data_out<= x"20";
        when x"2BE7" => data_out<= x"F0";
        when x"2BE8" => data_out<= x"80";
        when x"2BE9" => data_out<= x"A2";
        when x"2BEA" => data_out<= x"00";
        when x"2BEB" => data_out<= x"8A";
        when x"2BEC" => data_out<= x"20";
        when x"2BED" => data_out<= x"C3";
        when x"2BEE" => data_out<= x"B0";
        when x"2BEF" => data_out<= x"20";
        when x"2BF0" => data_out<= x"4C";
        when x"2BF1" => data_out<= x"AE";
        when x"2BF2" => data_out<= x"C9";
        when x"2BF3" => data_out<= x"50";
        when x"2BF4" => data_out<= x"8A";
        when x"2BF5" => data_out<= x"E9";
        when x"2BF6" => data_out<= x"C3";
        when x"2BF7" => data_out<= x"A5";
        when x"2BF8" => data_out<= x"0E";
        when x"2BF9" => data_out<= x"E9";
        when x"2BFA" => data_out<= x"00";
        when x"2BFB" => data_out<= x"A5";
        when x"2BFC" => data_out<= x"0F";
        when x"2BFD" => data_out<= x"E9";
        when x"2BFE" => data_out<= x"00";
        when x"2BFF" => data_out<= x"B0";
        when x"2C00" => data_out<= x"39";
        when x"2C01" => data_out<= x"20";
        when x"2C02" => data_out<= x"0A";
        when x"2C03" => data_out<= x"81";
        when x"2C04" => data_out<= x"AA";
        when x"2C05" => data_out<= x"F0";
        when x"2C06" => data_out<= x"26";
        when x"2C07" => data_out<= x"20";
        when x"2C08" => data_out<= x"FD";
        when x"2C09" => data_out<= x"80";
        when x"2C0A" => data_out<= x"A0";
        when x"2C0B" => data_out<= x"08";
        when x"2C0C" => data_out<= x"91";
        when x"2C0D" => data_out<= x"0C";
        when x"2C0E" => data_out<= x"C9";
        when x"2C0F" => data_out<= x"01";
        when x"2C10" => data_out<= x"F0";
        when x"2C11" => data_out<= x"38";
        when x"2C12" => data_out<= x"B1";
        when x"2C13" => data_out<= x"0C";
        when x"2C14" => data_out<= x"C9";
        when x"2C15" => data_out<= x"04";
        when x"2C16" => data_out<= x"D0";
        when x"2C17" => data_out<= x"08";
        when x"2C18" => data_out<= x"A9";
        when x"2C19" => data_out<= x"06";
        when x"2C1A" => data_out<= x"20";
        when x"2C1B" => data_out<= x"F0";
        when x"2C1C" => data_out<= x"80";
        when x"2C1D" => data_out<= x"4C";
        when x"2C1E" => data_out<= x"63";
        when x"2C1F" => data_out<= x"AD";
        when x"2C20" => data_out<= x"B1";
        when x"2C21" => data_out<= x"0C";
        when x"2C22" => data_out<= x"C9";
        when x"2C23" => data_out<= x"18";
        when x"2C24" => data_out<= x"D0";
        when x"2C25" => data_out<= x"07";
        when x"2C26" => data_out<= x"A2";
        when x"2C27" => data_out<= x"FF";
        when x"2C28" => data_out<= x"A9";
        when x"2C29" => data_out<= x"FE";
        when x"2C2A" => data_out<= x"4C";
        when x"2C2B" => data_out<= x"68";
        when x"2C2C" => data_out<= x"AD";
        when x"2C2D" => data_out<= x"20";
        when x"2C2E" => data_out<= x"4D";
        when x"2C2F" => data_out<= x"AF";
        when x"2C30" => data_out<= x"85";
        when x"2C31" => data_out<= x"10";
        when x"2C32" => data_out<= x"86";
        when x"2C33" => data_out<= x"11";
        when x"2C34" => data_out<= x"20";
        when x"2C35" => data_out<= x"E2";
        when x"2C36" => data_out<= x"AE";
        when x"2C37" => data_out<= x"4C";
        when x"2C38" => data_out<= x"EC";
        when x"2C39" => data_out<= x"AB";
        when x"2C3A" => data_out<= x"A0";
        when x"2C3B" => data_out<= x"02";
        when x"2C3C" => data_out<= x"B1";
        when x"2C3D" => data_out<= x"0C";
        when x"2C3E" => data_out<= x"18";
        when x"2C3F" => data_out<= x"69";
        when x"2C40" => data_out<= x"01";
        when x"2C41" => data_out<= x"4C";
        when x"2C42" => data_out<= x"DE";
        when x"2C43" => data_out<= x"AB";
        when x"2C44" => data_out<= x"A2";
        when x"2C45" => data_out<= x"FF";
        when x"2C46" => data_out<= x"8A";
        when x"2C47" => data_out<= x"4C";
        when x"2C48" => data_out<= x"68";
        when x"2C49" => data_out<= x"AD";
        when x"2C4A" => data_out<= x"20";
        when x"2C4B" => data_out<= x"FD";
        when x"2C4C" => data_out<= x"80";
        when x"2C4D" => data_out<= x"A0";
        when x"2C4E" => data_out<= x"07";
        when x"2C4F" => data_out<= x"91";
        when x"2C50" => data_out<= x"0C";
        when x"2C51" => data_out<= x"20";
        when x"2C52" => data_out<= x"FD";
        when x"2C53" => data_out<= x"80";
        when x"2C54" => data_out<= x"A0";
        when x"2C55" => data_out<= x"06";
        when x"2C56" => data_out<= x"91";
        when x"2C57" => data_out<= x"0C";
        when x"2C58" => data_out<= x"A9";
        when x"2C59" => data_out<= x"00";
        when x"2C5A" => data_out<= x"A0";
        when x"2C5B" => data_out<= x"04";
        when x"2C5C" => data_out<= x"91";
        when x"2C5D" => data_out<= x"0C";
        when x"2C5E" => data_out<= x"88";
        when x"2C5F" => data_out<= x"91";
        when x"2C60" => data_out<= x"0C";
        when x"2C61" => data_out<= x"C9";
        when x"2C62" => data_out<= x"80";
        when x"2C63" => data_out<= x"B0";
        when x"2C64" => data_out<= x"3A";
        when x"2C65" => data_out<= x"B1";
        when x"2C66" => data_out<= x"0C";
        when x"2C67" => data_out<= x"18";
        when x"2C68" => data_out<= x"A0";
        when x"2C69" => data_out<= x"0C";
        when x"2C6A" => data_out<= x"71";
        when x"2C6B" => data_out<= x"0C";
        when x"2C6C" => data_out<= x"48";
        when x"2C6D" => data_out<= x"A9";
        when x"2C6E" => data_out<= x"00";
        when x"2C6F" => data_out<= x"C8";
        when x"2C70" => data_out<= x"71";
        when x"2C71" => data_out<= x"0C";
        when x"2C72" => data_out<= x"AA";
        when x"2C73" => data_out<= x"68";
        when x"2C74" => data_out<= x"20";
        when x"2C75" => data_out<= x"7B";
        when x"2C76" => data_out<= x"B0";
        when x"2C77" => data_out<= x"20";
        when x"2C78" => data_out<= x"FD";
        when x"2C79" => data_out<= x"80";
        when x"2C7A" => data_out<= x"A0";
        when x"2C7B" => data_out<= x"00";
        when x"2C7C" => data_out<= x"20";
        when x"2C7D" => data_out<= x"AD";
        when x"2C7E" => data_out<= x"B0";
        when x"2C7F" => data_out<= x"A0";
        when x"2C80" => data_out<= x"0D";
        when x"2C81" => data_out<= x"20";
        when x"2C82" => data_out<= x"4F";
        when x"2C83" => data_out<= x"AF";
        when x"2C84" => data_out<= x"85";
        when x"2C85" => data_out<= x"14";
        when x"2C86" => data_out<= x"86";
        when x"2C87" => data_out<= x"15";
        when x"2C88" => data_out<= x"A0";
        when x"2C89" => data_out<= x"03";
        when x"2C8A" => data_out<= x"B1";
        when x"2C8B" => data_out<= x"0C";
        when x"2C8C" => data_out<= x"A8";
        when x"2C8D" => data_out<= x"B1";
        when x"2C8E" => data_out<= x"14";
        when x"2C8F" => data_out<= x"A0";
        when x"2C90" => data_out<= x"04";
        when x"2C91" => data_out<= x"18";
        when x"2C92" => data_out<= x"71";
        when x"2C93" => data_out<= x"0C";
        when x"2C94" => data_out<= x"91";
        when x"2C95" => data_out<= x"0C";
        when x"2C96" => data_out<= x"88";
        when x"2C97" => data_out<= x"B1";
        when x"2C98" => data_out<= x"0C";
        when x"2C99" => data_out<= x"18";
        when x"2C9A" => data_out<= x"69";
        when x"2C9B" => data_out<= x"01";
        when x"2C9C" => data_out<= x"4C";
        when x"2C9D" => data_out<= x"5F";
        when x"2C9E" => data_out<= x"AC";
        when x"2C9F" => data_out<= x"20";
        when x"2CA0" => data_out<= x"FD";
        when x"2CA1" => data_out<= x"80";
        when x"2CA2" => data_out<= x"A0";
        when x"2CA3" => data_out<= x"05";
        when x"2CA4" => data_out<= x"91";
        when x"2CA5" => data_out<= x"0C";
        when x"2CA6" => data_out<= x"A2";
        when x"2CA7" => data_out<= x"00";
        when x"2CA8" => data_out<= x"C8";
        when x"2CA9" => data_out<= x"B1";
        when x"2CAA" => data_out<= x"0C";
        when x"2CAB" => data_out<= x"18";
        when x"2CAC" => data_out<= x"C8";
        when x"2CAD" => data_out<= x"71";
        when x"2CAE" => data_out<= x"0C";
        when x"2CAF" => data_out<= x"90";
        when x"2CB0" => data_out<= x"01";
        when x"2CB1" => data_out<= x"E8";
        when x"2CB2" => data_out<= x"E0";
        when x"2CB3" => data_out<= x"00";
        when x"2CB4" => data_out<= x"D0";
        when x"2CB5" => data_out<= x"3E";
        when x"2CB6" => data_out<= x"C9";
        when x"2CB7" => data_out<= x"FF";
        when x"2CB8" => data_out<= x"D0";
        when x"2CB9" => data_out<= x"3A";
        when x"2CBA" => data_out<= x"A0";
        when x"2CBB" => data_out<= x"04";
        when x"2CBC" => data_out<= x"B1";
        when x"2CBD" => data_out<= x"0C";
        when x"2CBE" => data_out<= x"C8";
        when x"2CBF" => data_out<= x"D1";
        when x"2CC0" => data_out<= x"0C";
        when x"2CC1" => data_out<= x"D0";
        when x"2CC2" => data_out<= x"2F";
        when x"2CC3" => data_out<= x"A0";
        when x"2CC4" => data_out<= x"07";
        when x"2CC5" => data_out<= x"B1";
        when x"2CC6" => data_out<= x"0C";
        when x"2CC7" => data_out<= x"A0";
        when x"2CC8" => data_out<= x"0B";
        when x"2CC9" => data_out<= x"D1";
        when x"2CCA" => data_out<= x"0C";
        when x"2CCB" => data_out<= x"D0";
        when x"2CCC" => data_out<= x"25";
        when x"2CCD" => data_out<= x"A9";
        when x"2CCE" => data_out<= x"06";
        when x"2CCF" => data_out<= x"20";
        when x"2CD0" => data_out<= x"F0";
        when x"2CD1" => data_out<= x"80";
        when x"2CD2" => data_out<= x"A0";
        when x"2CD3" => data_out<= x"0C";
        when x"2CD4" => data_out<= x"A2";
        when x"2CD5" => data_out<= x"00";
        when x"2CD6" => data_out<= x"A9";
        when x"2CD7" => data_out<= x"80";
        when x"2CD8" => data_out<= x"20";
        when x"2CD9" => data_out<= x"04";
        when x"2CDA" => data_out<= x"AE";
        when x"2CDB" => data_out<= x"A0";
        when x"2CDC" => data_out<= x"09";
        when x"2CDD" => data_out<= x"A2";
        when x"2CDE" => data_out<= x"00";
        when x"2CDF" => data_out<= x"A9";
        when x"2CE0" => data_out<= x"80";
        when x"2CE1" => data_out<= x"20";
        when x"2CE2" => data_out<= x"04";
        when x"2CE3" => data_out<= x"AE";
        when x"2CE4" => data_out<= x"A0";
        when x"2CE5" => data_out<= x"0B";
        when x"2CE6" => data_out<= x"A2";
        when x"2CE7" => data_out<= x"00";
        when x"2CE8" => data_out<= x"B1";
        when x"2CE9" => data_out<= x"0C";
        when x"2CEA" => data_out<= x"18";
        when x"2CEB" => data_out<= x"69";
        when x"2CEC" => data_out<= x"01";
        when x"2CED" => data_out<= x"91";
        when x"2CEE" => data_out<= x"0C";
        when x"2CEF" => data_out<= x"4C";
        when x"2CF0" => data_out<= x"11";
        when x"2CF1" => data_out<= x"AD";
        when x"2CF2" => data_out<= x"A0";
        when x"2CF3" => data_out<= x"07";
        when x"2CF4" => data_out<= x"B1";
        when x"2CF5" => data_out<= x"0C";
        when x"2CF6" => data_out<= x"20";
        when x"2CF7" => data_out<= x"79";
        when x"2CF8" => data_out<= x"B0";
        when x"2CF9" => data_out<= x"A0";
        when x"2CFA" => data_out<= x"0D";
        when x"2CFB" => data_out<= x"B1";
        when x"2CFC" => data_out<= x"0C";
        when x"2CFD" => data_out<= x"38";
        when x"2CFE" => data_out<= x"E9";
        when x"2CFF" => data_out<= x"01";
        when x"2D00" => data_out<= x"20";
        when x"2D01" => data_out<= x"B4";
        when x"2D02" => data_out<= x"AE";
        when x"2D03" => data_out<= x"D0";
        when x"2D04" => data_out<= x"05";
        when x"2D05" => data_out<= x"A9";
        when x"2D06" => data_out<= x"06";
        when x"2D07" => data_out<= x"4C";
        when x"2D08" => data_out<= x"0C";
        when x"2D09" => data_out<= x"AD";
        when x"2D0A" => data_out<= x"A9";
        when x"2D0B" => data_out<= x"15";
        when x"2D0C" => data_out<= x"20";
        when x"2D0D" => data_out<= x"F0";
        when x"2D0E" => data_out<= x"80";
        when x"2D0F" => data_out<= x"A2";
        when x"2D10" => data_out<= x"00";
        when x"2D11" => data_out<= x"8A";
        when x"2D12" => data_out<= x"20";
        when x"2D13" => data_out<= x"C3";
        when x"2D14" => data_out<= x"B0";
        when x"2D15" => data_out<= x"20";
        when x"2D16" => data_out<= x"4C";
        when x"2D17" => data_out<= x"AE";
        when x"2D18" => data_out<= x"C9";
        when x"2D19" => data_out<= x"60";
        when x"2D1A" => data_out<= x"8A";
        when x"2D1B" => data_out<= x"E9";
        when x"2D1C" => data_out<= x"EA";
        when x"2D1D" => data_out<= x"A5";
        when x"2D1E" => data_out<= x"0E";
        when x"2D1F" => data_out<= x"E9";
        when x"2D20" => data_out<= x"00";
        when x"2D21" => data_out<= x"A5";
        when x"2D22" => data_out<= x"0F";
        when x"2D23" => data_out<= x"E9";
        when x"2D24" => data_out<= x"00";
        when x"2D25" => data_out<= x"B0";
        when x"2D26" => data_out<= x"3C";
        when x"2D27" => data_out<= x"20";
        when x"2D28" => data_out<= x"0A";
        when x"2D29" => data_out<= x"81";
        when x"2D2A" => data_out<= x"AA";
        when x"2D2B" => data_out<= x"F0";
        when x"2D2C" => data_out<= x"29";
        when x"2D2D" => data_out<= x"20";
        when x"2D2E" => data_out<= x"FD";
        when x"2D2F" => data_out<= x"80";
        when x"2D30" => data_out<= x"A0";
        when x"2D31" => data_out<= x"08";
        when x"2D32" => data_out<= x"91";
        when x"2D33" => data_out<= x"0C";
        when x"2D34" => data_out<= x"C9";
        when x"2D35" => data_out<= x"01";
        when x"2D36" => data_out<= x"D0";
        when x"2D37" => data_out<= x"03";
        when x"2D38" => data_out<= x"4C";
        when x"2D39" => data_out<= x"4A";
        when x"2D3A" => data_out<= x"AC";
        when x"2D3B" => data_out<= x"B1";
        when x"2D3C" => data_out<= x"0C";
        when x"2D3D" => data_out<= x"C9";
        when x"2D3E" => data_out<= x"04";
        when x"2D3F" => data_out<= x"D0";
        when x"2D40" => data_out<= x"08";
        when x"2D41" => data_out<= x"A9";
        when x"2D42" => data_out<= x"06";
        when x"2D43" => data_out<= x"20";
        when x"2D44" => data_out<= x"F0";
        when x"2D45" => data_out<= x"80";
        when x"2D46" => data_out<= x"4C";
        when x"2D47" => data_out<= x"63";
        when x"2D48" => data_out<= x"AD";
        when x"2D49" => data_out<= x"B1";
        when x"2D4A" => data_out<= x"0C";
        when x"2D4B" => data_out<= x"C9";
        when x"2D4C" => data_out<= x"18";
        when x"2D4D" => data_out<= x"D0";
        when x"2D4E" => data_out<= x"07";
        when x"2D4F" => data_out<= x"A2";
        when x"2D50" => data_out<= x"FF";
        when x"2D51" => data_out<= x"A9";
        when x"2D52" => data_out<= x"FE";
        when x"2D53" => data_out<= x"4C";
        when x"2D54" => data_out<= x"68";
        when x"2D55" => data_out<= x"AD";
        when x"2D56" => data_out<= x"20";
        when x"2D57" => data_out<= x"4D";
        when x"2D58" => data_out<= x"AF";
        when x"2D59" => data_out<= x"85";
        when x"2D5A" => data_out<= x"10";
        when x"2D5B" => data_out<= x"86";
        when x"2D5C" => data_out<= x"11";
        when x"2D5D" => data_out<= x"20";
        when x"2D5E" => data_out<= x"E2";
        when x"2D5F" => data_out<= x"AE";
        when x"2D60" => data_out<= x"4C";
        when x"2D61" => data_out<= x"12";
        when x"2D62" => data_out<= x"AD";
        when x"2D63" => data_out<= x"A0";
        when x"2D64" => data_out<= x"0A";
        when x"2D65" => data_out<= x"20";
        when x"2D66" => data_out<= x"4F";
        when x"2D67" => data_out<= x"AF";
        when x"2D68" => data_out<= x"A0";
        when x"2D69" => data_out<= x"10";
        when x"2D6A" => data_out<= x"4C";
        when x"2D6B" => data_out<= x"14";
        when x"2D6C" => data_out<= x"AE";
        when x"2D6D" => data_out<= x"A9";
        when x"2D6E" => data_out<= x"02";
        when x"2D6F" => data_out<= x"8D";
        when x"2D70" => data_out<= x"3C";
        when x"2D71" => data_out<= x"C0";
        when x"2D72" => data_out<= x"AD";
        when x"2D73" => data_out<= x"38";
        when x"2D74" => data_out<= x"C0";
        when x"2D75" => data_out<= x"AE";
        when x"2D76" => data_out<= x"39";
        when x"2D77" => data_out<= x"C0";
        when x"2D78" => data_out<= x"85";
        when x"2D79" => data_out<= x"0E";
        when x"2D7A" => data_out<= x"86";
        when x"2D7B" => data_out<= x"0F";
        when x"2D7C" => data_out<= x"AD";
        when x"2D7D" => data_out<= x"3A";
        when x"2D7E" => data_out<= x"C0";
        when x"2D7F" => data_out<= x"AE";
        when x"2D80" => data_out<= x"3B";
        when x"2D81" => data_out<= x"C0";
        when x"2D82" => data_out<= x"60";
        when x"2D83" => data_out<= x"85";
        when x"2D84" => data_out<= x"14";
        when x"2D85" => data_out<= x"86";
        when x"2D86" => data_out<= x"15";
        when x"2D87" => data_out<= x"20";
        when x"2D88" => data_out<= x"6D";
        when x"2D89" => data_out<= x"AD";
        when x"2D8A" => data_out<= x"18";
        when x"2D8B" => data_out<= x"65";
        when x"2D8C" => data_out<= x"14";
        when x"2D8D" => data_out<= x"85";
        when x"2D8E" => data_out<= x"08";
        when x"2D8F" => data_out<= x"8A";
        when x"2D90" => data_out<= x"65";
        when x"2D91" => data_out<= x"15";
        when x"2D92" => data_out<= x"85";
        when x"2D93" => data_out<= x"09";
        when x"2D94" => data_out<= x"A5";
        when x"2D95" => data_out<= x"0E";
        when x"2D96" => data_out<= x"69";
        when x"2D97" => data_out<= x"00";
        when x"2D98" => data_out<= x"85";
        when x"2D99" => data_out<= x"0A";
        when x"2D9A" => data_out<= x"A5";
        when x"2D9B" => data_out<= x"0F";
        when x"2D9C" => data_out<= x"69";
        when x"2D9D" => data_out<= x"00";
        when x"2D9E" => data_out<= x"85";
        when x"2D9F" => data_out<= x"0B";
        when x"2DA0" => data_out<= x"20";
        when x"2DA1" => data_out<= x"6D";
        when x"2DA2" => data_out<= x"AD";
        when x"2DA3" => data_out<= x"85";
        when x"2DA4" => data_out<= x"14";
        when x"2DA5" => data_out<= x"86";
        when x"2DA6" => data_out<= x"15";
        when x"2DA7" => data_out<= x"A5";
        when x"2DA8" => data_out<= x"0F";
        when x"2DA9" => data_out<= x"C5";
        when x"2DAA" => data_out<= x"0B";
        when x"2DAB" => data_out<= x"90";
        when x"2DAC" => data_out<= x"F3";
        when x"2DAD" => data_out<= x"D0";
        when x"2DAE" => data_out<= x"16";
        when x"2DAF" => data_out<= x"A5";
        when x"2DB0" => data_out<= x"0E";
        when x"2DB1" => data_out<= x"C5";
        when x"2DB2" => data_out<= x"0A";
        when x"2DB3" => data_out<= x"90";
        when x"2DB4" => data_out<= x"EB";
        when x"2DB5" => data_out<= x"D0";
        when x"2DB6" => data_out<= x"0E";
        when x"2DB7" => data_out<= x"A5";
        when x"2DB8" => data_out<= x"15";
        when x"2DB9" => data_out<= x"C5";
        when x"2DBA" => data_out<= x"09";
        when x"2DBB" => data_out<= x"90";
        when x"2DBC" => data_out<= x"E3";
        when x"2DBD" => data_out<= x"D0";
        when x"2DBE" => data_out<= x"06";
        when x"2DBF" => data_out<= x"A5";
        when x"2DC0" => data_out<= x"14";
        when x"2DC1" => data_out<= x"C5";
        when x"2DC2" => data_out<= x"08";
        when x"2DC3" => data_out<= x"90";
        when x"2DC4" => data_out<= x"DB";
        when x"2DC5" => data_out<= x"60";
        when x"2DC6" => data_out<= x"85";
        when x"2DC7" => data_out<= x"14";
        when x"2DC8" => data_out<= x"86";
        when x"2DC9" => data_out<= x"15";
        when x"2DCA" => data_out<= x"05";
        when x"2DCB" => data_out<= x"15";
        when x"2DCC" => data_out<= x"F0";
        when x"2DCD" => data_out<= x"15";
        when x"2DCE" => data_out<= x"A9";
        when x"2DCF" => data_out<= x"E8";
        when x"2DD0" => data_out<= x"A2";
        when x"2DD1" => data_out<= x"03";
        when x"2DD2" => data_out<= x"20";
        when x"2DD3" => data_out<= x"83";
        when x"2DD4" => data_out<= x"AD";
        when x"2DD5" => data_out<= x"A5";
        when x"2DD6" => data_out<= x"14";
        when x"2DD7" => data_out<= x"D0";
        when x"2DD8" => data_out<= x"02";
        when x"2DD9" => data_out<= x"C6";
        when x"2DDA" => data_out<= x"15";
        when x"2DDB" => data_out<= x"C6";
        when x"2DDC" => data_out<= x"14";
        when x"2DDD" => data_out<= x"A5";
        when x"2DDE" => data_out<= x"14";
        when x"2DDF" => data_out<= x"05";
        when x"2DE0" => data_out<= x"15";
        when x"2DE1" => data_out<= x"D0";
        when x"2DE2" => data_out<= x"EB";
        when x"2DE3" => data_out<= x"60";
        when x"2DE4" => data_out<= x"40";
        when x"2DE5" => data_out<= x"40";
        when x"2DE6" => data_out<= x"A2";
        when x"2DE7" => data_out<= x"00";
        when x"2DE8" => data_out<= x"18";
        when x"2DE9" => data_out<= x"A0";
        when x"2DEA" => data_out<= x"00";
        when x"2DEB" => data_out<= x"71";
        when x"2DEC" => data_out<= x"0C";
        when x"2DED" => data_out<= x"C8";
        when x"2DEE" => data_out<= x"85";
        when x"2DEF" => data_out<= x"1C";
        when x"2DF0" => data_out<= x"8A";
        when x"2DF1" => data_out<= x"71";
        when x"2DF2" => data_out<= x"0C";
        when x"2DF3" => data_out<= x"AA";
        when x"2DF4" => data_out<= x"18";
        when x"2DF5" => data_out<= x"A5";
        when x"2DF6" => data_out<= x"0C";
        when x"2DF7" => data_out<= x"69";
        when x"2DF8" => data_out<= x"02";
        when x"2DF9" => data_out<= x"85";
        when x"2DFA" => data_out<= x"0C";
        when x"2DFB" => data_out<= x"90";
        when x"2DFC" => data_out<= x"02";
        when x"2DFD" => data_out<= x"E6";
        when x"2DFE" => data_out<= x"0D";
        when x"2DFF" => data_out<= x"A5";
        when x"2E00" => data_out<= x"1C";
        when x"2E01" => data_out<= x"60";
        when x"2E02" => data_out<= x"A0";
        when x"2E03" => data_out<= x"00";
        when x"2E04" => data_out<= x"18";
        when x"2E05" => data_out<= x"71";
        when x"2E06" => data_out<= x"0C";
        when x"2E07" => data_out<= x"91";
        when x"2E08" => data_out<= x"0C";
        when x"2E09" => data_out<= x"48";
        when x"2E0A" => data_out<= x"C8";
        when x"2E0B" => data_out<= x"8A";
        when x"2E0C" => data_out<= x"71";
        when x"2E0D" => data_out<= x"0C";
        when x"2E0E" => data_out<= x"91";
        when x"2E0F" => data_out<= x"0C";
        when x"2E10" => data_out<= x"AA";
        when x"2E11" => data_out<= x"68";
        when x"2E12" => data_out<= x"60";
        when x"2E13" => data_out<= x"C8";
        when x"2E14" => data_out<= x"48";
        when x"2E15" => data_out<= x"18";
        when x"2E16" => data_out<= x"98";
        when x"2E17" => data_out<= x"65";
        when x"2E18" => data_out<= x"0C";
        when x"2E19" => data_out<= x"85";
        when x"2E1A" => data_out<= x"0C";
        when x"2E1B" => data_out<= x"90";
        when x"2E1C" => data_out<= x"02";
        when x"2E1D" => data_out<= x"E6";
        when x"2E1E" => data_out<= x"0D";
        when x"2E1F" => data_out<= x"68";
        when x"2E20" => data_out<= x"60";
        when x"2E21" => data_out<= x"86";
        when x"2E22" => data_out<= x"1C";
        when x"2E23" => data_out<= x"0A";
        when x"2E24" => data_out<= x"26";
        when x"2E25" => data_out<= x"1C";
        when x"2E26" => data_out<= x"A6";
        when x"2E27" => data_out<= x"1C";
        when x"2E28" => data_out<= x"60";
        when x"2E29" => data_out<= x"86";
        when x"2E2A" => data_out<= x"1C";
        when x"2E2B" => data_out<= x"0A";
        when x"2E2C" => data_out<= x"26";
        when x"2E2D" => data_out<= x"1C";
        when x"2E2E" => data_out<= x"0A";
        when x"2E2F" => data_out<= x"26";
        when x"2E30" => data_out<= x"1C";
        when x"2E31" => data_out<= x"0A";
        when x"2E32" => data_out<= x"26";
        when x"2E33" => data_out<= x"1C";
        when x"2E34" => data_out<= x"0A";
        when x"2E35" => data_out<= x"26";
        when x"2E36" => data_out<= x"1C";
        when x"2E37" => data_out<= x"A6";
        when x"2E38" => data_out<= x"1C";
        when x"2E39" => data_out<= x"60";
        when x"2E3A" => data_out<= x"86";
        when x"2E3B" => data_out<= x"1C";
        when x"2E3C" => data_out<= x"0A";
        when x"2E3D" => data_out<= x"26";
        when x"2E3E" => data_out<= x"1C";
        when x"2E3F" => data_out<= x"26";
        when x"2E40" => data_out<= x"0E";
        when x"2E41" => data_out<= x"26";
        when x"2E42" => data_out<= x"0F";
        when x"2E43" => data_out<= x"A6";
        when x"2E44" => data_out<= x"1C";
        when x"2E45" => data_out<= x"60";
        when x"2E46" => data_out<= x"A0";
        when x"2E47" => data_out<= x"FF";
        when x"2E48" => data_out<= x"E0";
        when x"2E49" => data_out<= x"80";
        when x"2E4A" => data_out<= x"B0";
        when x"2E4B" => data_out<= x"02";
        when x"2E4C" => data_out<= x"A0";
        when x"2E4D" => data_out<= x"00";
        when x"2E4E" => data_out<= x"84";
        when x"2E4F" => data_out<= x"0E";
        when x"2E50" => data_out<= x"84";
        when x"2E51" => data_out<= x"0F";
        when x"2E52" => data_out<= x"60";
        when x"2E53" => data_out<= x"85";
        when x"2E54" => data_out<= x"14";
        when x"2E55" => data_out<= x"86";
        when x"2E56" => data_out<= x"15";
        when x"2E57" => data_out<= x"6C";
        when x"2E58" => data_out<= x"14";
        when x"2E59" => data_out<= x"00";
        when x"2E5A" => data_out<= x"38";
        when x"2E5B" => data_out<= x"E9";
        when x"2E5C" => data_out<= x"01";
        when x"2E5D" => data_out<= x"B0";
        when x"2E5E" => data_out<= x"01";
        when x"2E5F" => data_out<= x"CA";
        when x"2E60" => data_out<= x"60";
        when x"2E61" => data_out<= x"84";
        when x"2E62" => data_out<= x"1C";
        when x"2E63" => data_out<= x"38";
        when x"2E64" => data_out<= x"E5";
        when x"2E65" => data_out<= x"1C";
        when x"2E66" => data_out<= x"B0";
        when x"2E67" => data_out<= x"01";
        when x"2E68" => data_out<= x"CA";
        when x"2E69" => data_out<= x"60";
        when x"2E6A" => data_out<= x"A4";
        when x"2E6B" => data_out<= x"0C";
        when x"2E6C" => data_out<= x"D0";
        when x"2E6D" => data_out<= x"02";
        when x"2E6E" => data_out<= x"C6";
        when x"2E6F" => data_out<= x"0D";
        when x"2E70" => data_out<= x"C6";
        when x"2E71" => data_out<= x"0C";
        when x"2E72" => data_out<= x"60";
        when x"2E73" => data_out<= x"A5";
        when x"2E74" => data_out<= x"0C";
        when x"2E75" => data_out<= x"38";
        when x"2E76" => data_out<= x"E9";
        when x"2E77" => data_out<= x"02";
        when x"2E78" => data_out<= x"85";
        when x"2E79" => data_out<= x"0C";
        when x"2E7A" => data_out<= x"90";
        when x"2E7B" => data_out<= x"01";
        when x"2E7C" => data_out<= x"60";
        when x"2E7D" => data_out<= x"C6";
        when x"2E7E" => data_out<= x"0D";
        when x"2E7F" => data_out<= x"60";
        when x"2E80" => data_out<= x"A5";
        when x"2E81" => data_out<= x"0C";
        when x"2E82" => data_out<= x"38";
        when x"2E83" => data_out<= x"E9";
        when x"2E84" => data_out<= x"03";
        when x"2E85" => data_out<= x"85";
        when x"2E86" => data_out<= x"0C";
        when x"2E87" => data_out<= x"90";
        when x"2E88" => data_out<= x"01";
        when x"2E89" => data_out<= x"60";
        when x"2E8A" => data_out<= x"C6";
        when x"2E8B" => data_out<= x"0D";
        when x"2E8C" => data_out<= x"60";
        when x"2E8D" => data_out<= x"A5";
        when x"2E8E" => data_out<= x"0C";
        when x"2E8F" => data_out<= x"38";
        when x"2E90" => data_out<= x"E9";
        when x"2E91" => data_out<= x"04";
        when x"2E92" => data_out<= x"85";
        when x"2E93" => data_out<= x"0C";
        when x"2E94" => data_out<= x"90";
        when x"2E95" => data_out<= x"01";
        when x"2E96" => data_out<= x"60";
        when x"2E97" => data_out<= x"C6";
        when x"2E98" => data_out<= x"0D";
        when x"2E99" => data_out<= x"60";
        when x"2E9A" => data_out<= x"A5";
        when x"2E9B" => data_out<= x"0C";
        when x"2E9C" => data_out<= x"38";
        when x"2E9D" => data_out<= x"E9";
        when x"2E9E" => data_out<= x"06";
        when x"2E9F" => data_out<= x"85";
        when x"2EA0" => data_out<= x"0C";
        when x"2EA1" => data_out<= x"90";
        when x"2EA2" => data_out<= x"01";
        when x"2EA3" => data_out<= x"60";
        when x"2EA4" => data_out<= x"C6";
        when x"2EA5" => data_out<= x"0D";
        when x"2EA6" => data_out<= x"60";
        when x"2EA7" => data_out<= x"A5";
        when x"2EA8" => data_out<= x"0C";
        when x"2EA9" => data_out<= x"38";
        when x"2EAA" => data_out<= x"E9";
        when x"2EAB" => data_out<= x"07";
        when x"2EAC" => data_out<= x"85";
        when x"2EAD" => data_out<= x"0C";
        when x"2EAE" => data_out<= x"90";
        when x"2EAF" => data_out<= x"01";
        when x"2EB0" => data_out<= x"60";
        when x"2EB1" => data_out<= x"C6";
        when x"2EB2" => data_out<= x"0D";
        when x"2EB3" => data_out<= x"60";
        when x"2EB4" => data_out<= x"A2";
        when x"2EB5" => data_out<= x"00";
        when x"2EB6" => data_out<= x"85";
        when x"2EB7" => data_out<= x"0E";
        when x"2EB8" => data_out<= x"86";
        when x"2EB9" => data_out<= x"0F";
        when x"2EBA" => data_out<= x"A0";
        when x"2EBB" => data_out<= x"00";
        when x"2EBC" => data_out<= x"B1";
        when x"2EBD" => data_out<= x"0C";
        when x"2EBE" => data_out<= x"AA";
        when x"2EBF" => data_out<= x"E6";
        when x"2EC0" => data_out<= x"0C";
        when x"2EC1" => data_out<= x"D0";
        when x"2EC2" => data_out<= x"02";
        when x"2EC3" => data_out<= x"E6";
        when x"2EC4" => data_out<= x"0D";
        when x"2EC5" => data_out<= x"B1";
        when x"2EC6" => data_out<= x"0C";
        when x"2EC7" => data_out<= x"E6";
        when x"2EC8" => data_out<= x"0C";
        when x"2EC9" => data_out<= x"D0";
        when x"2ECA" => data_out<= x"02";
        when x"2ECB" => data_out<= x"E6";
        when x"2ECC" => data_out<= x"0D";
        when x"2ECD" => data_out<= x"38";
        when x"2ECE" => data_out<= x"E5";
        when x"2ECF" => data_out<= x"0F";
        when x"2ED0" => data_out<= x"D0";
        when x"2ED1" => data_out<= x"09";
        when x"2ED2" => data_out<= x"E4";
        when x"2ED3" => data_out<= x"0E";
        when x"2ED4" => data_out<= x"F0";
        when x"2ED5" => data_out<= x"04";
        when x"2ED6" => data_out<= x"69";
        when x"2ED7" => data_out<= x"FF";
        when x"2ED8" => data_out<= x"09";
        when x"2ED9" => data_out<= x"01";
        when x"2EDA" => data_out<= x"60";
        when x"2EDB" => data_out<= x"50";
        when x"2EDC" => data_out<= x"FD";
        when x"2EDD" => data_out<= x"49";
        when x"2EDE" => data_out<= x"FF";
        when x"2EDF" => data_out<= x"09";
        when x"2EE0" => data_out<= x"01";
        when x"2EE1" => data_out<= x"60";
        when x"2EE2" => data_out<= x"18";
        when x"2EE3" => data_out<= x"69";
        when x"2EE4" => data_out<= x"01";
        when x"2EE5" => data_out<= x"90";
        when x"2EE6" => data_out<= x"01";
        when x"2EE7" => data_out<= x"E8";
        when x"2EE8" => data_out<= x"60";
        when x"2EE9" => data_out<= x"18";
        when x"2EEA" => data_out<= x"69";
        when x"2EEB" => data_out<= x"02";
        when x"2EEC" => data_out<= x"90";
        when x"2EED" => data_out<= x"01";
        when x"2EEE" => data_out<= x"E8";
        when x"2EEF" => data_out<= x"60";
        when x"2EF0" => data_out<= x"A0";
        when x"2EF1" => data_out<= x"03";
        when x"2EF2" => data_out<= x"4C";
        when x"2EF3" => data_out<= x"FC";
        when x"2EF4" => data_out<= x"AE";
        when x"2EF5" => data_out<= x"A0";
        when x"2EF6" => data_out<= x"05";
        when x"2EF7" => data_out<= x"4C";
        when x"2EF8" => data_out<= x"FC";
        when x"2EF9" => data_out<= x"AE";
        when x"2EFA" => data_out<= x"A0";
        when x"2EFB" => data_out<= x"04";
        when x"2EFC" => data_out<= x"84";
        when x"2EFD" => data_out<= x"1C";
        when x"2EFE" => data_out<= x"18";
        when x"2EFF" => data_out<= x"65";
        when x"2F00" => data_out<= x"1C";
        when x"2F01" => data_out<= x"90";
        when x"2F02" => data_out<= x"01";
        when x"2F03" => data_out<= x"E8";
        when x"2F04" => data_out<= x"60";
        when x"2F05" => data_out<= x"E6";
        when x"2F06" => data_out<= x"0C";
        when x"2F07" => data_out<= x"D0";
        when x"2F08" => data_out<= x"02";
        when x"2F09" => data_out<= x"E6";
        when x"2F0A" => data_out<= x"0D";
        when x"2F0B" => data_out<= x"60";
        when x"2F0C" => data_out<= x"A0";
        when x"2F0D" => data_out<= x"01";
        when x"2F0E" => data_out<= x"B1";
        when x"2F0F" => data_out<= x"0C";
        when x"2F10" => data_out<= x"AA";
        when x"2F11" => data_out<= x"88";
        when x"2F12" => data_out<= x"B1";
        when x"2F13" => data_out<= x"0C";
        when x"2F14" => data_out<= x"E6";
        when x"2F15" => data_out<= x"0C";
        when x"2F16" => data_out<= x"F0";
        when x"2F17" => data_out<= x"05";
        when x"2F18" => data_out<= x"E6";
        when x"2F19" => data_out<= x"0C";
        when x"2F1A" => data_out<= x"F0";
        when x"2F1B" => data_out<= x"03";
        when x"2F1C" => data_out<= x"60";
        when x"2F1D" => data_out<= x"E6";
        when x"2F1E" => data_out<= x"0C";
        when x"2F1F" => data_out<= x"E6";
        when x"2F20" => data_out<= x"0D";
        when x"2F21" => data_out<= x"60";
        when x"2F22" => data_out<= x"A0";
        when x"2F23" => data_out<= x"03";
        when x"2F24" => data_out<= x"4C";
        when x"2F25" => data_out<= x"14";
        when x"2F26" => data_out<= x"AE";
        when x"2F27" => data_out<= x"A0";
        when x"2F28" => data_out<= x"04";
        when x"2F29" => data_out<= x"4C";
        when x"2F2A" => data_out<= x"14";
        when x"2F2B" => data_out<= x"AE";
        when x"2F2C" => data_out<= x"A0";
        when x"2F2D" => data_out<= x"05";
        when x"2F2E" => data_out<= x"4C";
        when x"2F2F" => data_out<= x"14";
        when x"2F30" => data_out<= x"AE";
        when x"2F31" => data_out<= x"A0";
        when x"2F32" => data_out<= x"06";
        when x"2F33" => data_out<= x"4C";
        when x"2F34" => data_out<= x"14";
        when x"2F35" => data_out<= x"AE";
        when x"2F36" => data_out<= x"A0";
        when x"2F37" => data_out<= x"07";
        when x"2F38" => data_out<= x"4C";
        when x"2F39" => data_out<= x"14";
        when x"2F3A" => data_out<= x"AE";
        when x"2F3B" => data_out<= x"A0";
        when x"2F3C" => data_out<= x"08";
        when x"2F3D" => data_out<= x"4C";
        when x"2F3E" => data_out<= x"14";
        when x"2F3F" => data_out<= x"AE";
        when x"2F40" => data_out<= x"A0";
        when x"2F41" => data_out<= x"01";
        when x"2F42" => data_out<= x"85";
        when x"2F43" => data_out<= x"14";
        when x"2F44" => data_out<= x"86";
        when x"2F45" => data_out<= x"15";
        when x"2F46" => data_out<= x"B1";
        when x"2F47" => data_out<= x"14";
        when x"2F48" => data_out<= x"AA";
        when x"2F49" => data_out<= x"88";
        when x"2F4A" => data_out<= x"B1";
        when x"2F4B" => data_out<= x"14";
        when x"2F4C" => data_out<= x"60";
        when x"2F4D" => data_out<= x"A0";
        when x"2F4E" => data_out<= x"01";
        when x"2F4F" => data_out<= x"B1";
        when x"2F50" => data_out<= x"0C";
        when x"2F51" => data_out<= x"AA";
        when x"2F52" => data_out<= x"88";
        when x"2F53" => data_out<= x"B1";
        when x"2F54" => data_out<= x"0C";
        when x"2F55" => data_out<= x"60";
        when x"2F56" => data_out<= x"A0";
        when x"2F57" => data_out<= x"03";
        when x"2F58" => data_out<= x"B1";
        when x"2F59" => data_out<= x"0C";
        when x"2F5A" => data_out<= x"85";
        when x"2F5B" => data_out<= x"0F";
        when x"2F5C" => data_out<= x"88";
        when x"2F5D" => data_out<= x"B1";
        when x"2F5E" => data_out<= x"0C";
        when x"2F5F" => data_out<= x"85";
        when x"2F60" => data_out<= x"0E";
        when x"2F61" => data_out<= x"88";
        when x"2F62" => data_out<= x"B1";
        when x"2F63" => data_out<= x"0C";
        when x"2F64" => data_out<= x"AA";
        when x"2F65" => data_out<= x"88";
        when x"2F66" => data_out<= x"B1";
        when x"2F67" => data_out<= x"0C";
        when x"2F68" => data_out<= x"60";
        when x"2F69" => data_out<= x"A2";
        when x"2F6A" => data_out<= x"00";
        when x"2F6B" => data_out<= x"18";
        when x"2F6C" => data_out<= x"65";
        when x"2F6D" => data_out<= x"0C";
        when x"2F6E" => data_out<= x"48";
        when x"2F6F" => data_out<= x"8A";
        when x"2F70" => data_out<= x"65";
        when x"2F71" => data_out<= x"0D";
        when x"2F72" => data_out<= x"AA";
        when x"2F73" => data_out<= x"68";
        when x"2F74" => data_out<= x"60";
        when x"2F75" => data_out<= x"A9";
        when x"2F76" => data_out<= x"00";
        when x"2F77" => data_out<= x"AA";
        when x"2F78" => data_out<= x"A0";
        when x"2F79" => data_out<= x"00";
        when x"2F7A" => data_out<= x"84";
        when x"2F7B" => data_out<= x"0E";
        when x"2F7C" => data_out<= x"84";
        when x"2F7D" => data_out<= x"0F";
        when x"2F7E" => data_out<= x"48";
        when x"2F7F" => data_out<= x"20";
        when x"2F80" => data_out<= x"8D";
        when x"2F81" => data_out<= x"AE";
        when x"2F82" => data_out<= x"A0";
        when x"2F83" => data_out<= x"03";
        when x"2F84" => data_out<= x"A5";
        when x"2F85" => data_out<= x"0F";
        when x"2F86" => data_out<= x"91";
        when x"2F87" => data_out<= x"0C";
        when x"2F88" => data_out<= x"88";
        when x"2F89" => data_out<= x"A5";
        when x"2F8A" => data_out<= x"0E";
        when x"2F8B" => data_out<= x"91";
        when x"2F8C" => data_out<= x"0C";
        when x"2F8D" => data_out<= x"88";
        when x"2F8E" => data_out<= x"8A";
        when x"2F8F" => data_out<= x"91";
        when x"2F90" => data_out<= x"0C";
        when x"2F91" => data_out<= x"68";
        when x"2F92" => data_out<= x"88";
        when x"2F93" => data_out<= x"91";
        when x"2F94" => data_out<= x"0C";
        when x"2F95" => data_out<= x"60";
        when x"2F96" => data_out<= x"20";
        when x"2F97" => data_out<= x"BF";
        when x"2F98" => data_out<= x"AF";
        when x"2F99" => data_out<= x"A6";
        when x"2F9A" => data_out<= x"19";
        when x"2F9B" => data_out<= x"F0";
        when x"2F9C" => data_out<= x"13";
        when x"2F9D" => data_out<= x"B1";
        when x"2F9E" => data_out<= x"14";
        when x"2F9F" => data_out<= x"91";
        when x"2FA0" => data_out<= x"16";
        when x"2FA1" => data_out<= x"C8";
        when x"2FA2" => data_out<= x"B1";
        when x"2FA3" => data_out<= x"14";
        when x"2FA4" => data_out<= x"91";
        when x"2FA5" => data_out<= x"16";
        when x"2FA6" => data_out<= x"C8";
        when x"2FA7" => data_out<= x"D0";
        when x"2FA8" => data_out<= x"F4";
        when x"2FA9" => data_out<= x"E6";
        when x"2FAA" => data_out<= x"15";
        when x"2FAB" => data_out<= x"E6";
        when x"2FAC" => data_out<= x"17";
        when x"2FAD" => data_out<= x"CA";
        when x"2FAE" => data_out<= x"D0";
        when x"2FAF" => data_out<= x"ED";
        when x"2FB0" => data_out<= x"A6";
        when x"2FB1" => data_out<= x"18";
        when x"2FB2" => data_out<= x"F0";
        when x"2FB3" => data_out<= x"08";
        when x"2FB4" => data_out<= x"B1";
        when x"2FB5" => data_out<= x"14";
        when x"2FB6" => data_out<= x"91";
        when x"2FB7" => data_out<= x"16";
        when x"2FB8" => data_out<= x"C8";
        when x"2FB9" => data_out<= x"CA";
        when x"2FBA" => data_out<= x"D0";
        when x"2FBB" => data_out<= x"F8";
        when x"2FBC" => data_out<= x"4C";
        when x"2FBD" => data_out<= x"0C";
        when x"2FBE" => data_out<= x"AF";
        when x"2FBF" => data_out<= x"85";
        when x"2FC0" => data_out<= x"18";
        when x"2FC1" => data_out<= x"86";
        when x"2FC2" => data_out<= x"19";
        when x"2FC3" => data_out<= x"20";
        when x"2FC4" => data_out<= x"53";
        when x"2FC5" => data_out<= x"B0";
        when x"2FC6" => data_out<= x"C8";
        when x"2FC7" => data_out<= x"B1";
        when x"2FC8" => data_out<= x"0C";
        when x"2FC9" => data_out<= x"AA";
        when x"2FCA" => data_out<= x"86";
        when x"2FCB" => data_out<= x"17";
        when x"2FCC" => data_out<= x"88";
        when x"2FCD" => data_out<= x"B1";
        when x"2FCE" => data_out<= x"0C";
        when x"2FCF" => data_out<= x"85";
        when x"2FD0" => data_out<= x"16";
        when x"2FD1" => data_out<= x"60";
        when x"2FD2" => data_out<= x"85";
        when x"2FD3" => data_out<= x"18";
        when x"2FD4" => data_out<= x"86";
        when x"2FD5" => data_out<= x"19";
        when x"2FD6" => data_out<= x"A2";
        when x"2FD7" => data_out<= x"00";
        when x"2FD8" => data_out<= x"F0";
        when x"2FD9" => data_out<= x"08";
        when x"2FDA" => data_out<= x"85";
        when x"2FDB" => data_out<= x"18";
        when x"2FDC" => data_out<= x"86";
        when x"2FDD" => data_out<= x"19";
        when x"2FDE" => data_out<= x"20";
        when x"2FDF" => data_out<= x"0C";
        when x"2FE0" => data_out<= x"AF";
        when x"2FE1" => data_out<= x"AA";
        when x"2FE2" => data_out<= x"A0";
        when x"2FE3" => data_out<= x"01";
        when x"2FE4" => data_out<= x"B1";
        when x"2FE5" => data_out<= x"0C";
        when x"2FE6" => data_out<= x"85";
        when x"2FE7" => data_out<= x"15";
        when x"2FE8" => data_out<= x"88";
        when x"2FE9" => data_out<= x"B1";
        when x"2FEA" => data_out<= x"0C";
        when x"2FEB" => data_out<= x"85";
        when x"2FEC" => data_out<= x"14";
        when x"2FED" => data_out<= x"46";
        when x"2FEE" => data_out<= x"19";
        when x"2FEF" => data_out<= x"66";
        when x"2FF0" => data_out<= x"18";
        when x"2FF1" => data_out<= x"90";
        when x"2FF2" => data_out<= x"09";
        when x"2FF3" => data_out<= x"8A";
        when x"2FF4" => data_out<= x"91";
        when x"2FF5" => data_out<= x"14";
        when x"2FF6" => data_out<= x"E6";
        when x"2FF7" => data_out<= x"14";
        when x"2FF8" => data_out<= x"D0";
        when x"2FF9" => data_out<= x"02";
        when x"2FFA" => data_out<= x"E6";
        when x"2FFB" => data_out<= x"15";
        when x"2FFC" => data_out<= x"A5";
        when x"2FFD" => data_out<= x"14";
        when x"2FFE" => data_out<= x"18";
        when x"2FFF" => data_out<= x"65";
        when x"3000" => data_out<= x"18";
        when x"3001" => data_out<= x"85";
        when x"3002" => data_out<= x"16";
        when x"3003" => data_out<= x"A5";
        when x"3004" => data_out<= x"15";
        when x"3005" => data_out<= x"65";
        when x"3006" => data_out<= x"19";
        when x"3007" => data_out<= x"85";
        when x"3008" => data_out<= x"17";
        when x"3009" => data_out<= x"8A";
        when x"300A" => data_out<= x"A6";
        when x"300B" => data_out<= x"19";
        when x"300C" => data_out<= x"F0";
        when x"300D" => data_out<= x"13";
        when x"300E" => data_out<= x"91";
        when x"300F" => data_out<= x"14";
        when x"3010" => data_out<= x"91";
        when x"3011" => data_out<= x"16";
        when x"3012" => data_out<= x"C8";
        when x"3013" => data_out<= x"91";
        when x"3014" => data_out<= x"14";
        when x"3015" => data_out<= x"91";
        when x"3016" => data_out<= x"16";
        when x"3017" => data_out<= x"C8";
        when x"3018" => data_out<= x"D0";
        when x"3019" => data_out<= x"F4";
        when x"301A" => data_out<= x"E6";
        when x"301B" => data_out<= x"15";
        when x"301C" => data_out<= x"E6";
        when x"301D" => data_out<= x"17";
        when x"301E" => data_out<= x"CA";
        when x"301F" => data_out<= x"D0";
        when x"3020" => data_out<= x"ED";
        when x"3021" => data_out<= x"A4";
        when x"3022" => data_out<= x"18";
        when x"3023" => data_out<= x"F0";
        when x"3024" => data_out<= x"07";
        when x"3025" => data_out<= x"88";
        when x"3026" => data_out<= x"91";
        when x"3027" => data_out<= x"14";
        when x"3028" => data_out<= x"91";
        when x"3029" => data_out<= x"16";
        when x"302A" => data_out<= x"D0";
        when x"302B" => data_out<= x"F9";
        when x"302C" => data_out<= x"4C";
        when x"302D" => data_out<= x"0C";
        when x"302E" => data_out<= x"AF";
        when x"302F" => data_out<= x"E0";
        when x"3030" => data_out<= x"00";
        when x"3031" => data_out<= x"10";
        when x"3032" => data_out<= x"0D";
        when x"3033" => data_out<= x"18";
        when x"3034" => data_out<= x"49";
        when x"3035" => data_out<= x"FF";
        when x"3036" => data_out<= x"69";
        when x"3037" => data_out<= x"01";
        when x"3038" => data_out<= x"48";
        when x"3039" => data_out<= x"8A";
        when x"303A" => data_out<= x"49";
        when x"303B" => data_out<= x"FF";
        when x"303C" => data_out<= x"69";
        when x"303D" => data_out<= x"00";
        when x"303E" => data_out<= x"AA";
        when x"303F" => data_out<= x"68";
        when x"3040" => data_out<= x"60";
        when x"3041" => data_out<= x"A2";
        when x"3042" => data_out<= x"00";
        when x"3043" => data_out<= x"A0";
        when x"3044" => data_out<= x"00";
        when x"3045" => data_out<= x"11";
        when x"3046" => data_out<= x"0C";
        when x"3047" => data_out<= x"C8";
        when x"3048" => data_out<= x"85";
        when x"3049" => data_out<= x"1C";
        when x"304A" => data_out<= x"8A";
        when x"304B" => data_out<= x"11";
        when x"304C" => data_out<= x"0C";
        when x"304D" => data_out<= x"AA";
        when x"304E" => data_out<= x"A5";
        when x"304F" => data_out<= x"1C";
        when x"3050" => data_out<= x"4C";
        when x"3051" => data_out<= x"13";
        when x"3052" => data_out<= x"AE";
        when x"3053" => data_out<= x"A0";
        when x"3054" => data_out<= x"01";
        when x"3055" => data_out<= x"B1";
        when x"3056" => data_out<= x"0C";
        when x"3057" => data_out<= x"85";
        when x"3058" => data_out<= x"15";
        when x"3059" => data_out<= x"88";
        when x"305A" => data_out<= x"B1";
        when x"305B" => data_out<= x"0C";
        when x"305C" => data_out<= x"85";
        when x"305D" => data_out<= x"14";
        when x"305E" => data_out<= x"4C";
        when x"305F" => data_out<= x"14";
        when x"3060" => data_out<= x"AF";
        when x"3061" => data_out<= x"A0";
        when x"3062" => data_out<= x"00";
        when x"3063" => data_out<= x"B1";
        when x"3064" => data_out<= x"0C";
        when x"3065" => data_out<= x"A4";
        when x"3066" => data_out<= x"0C";
        when x"3067" => data_out<= x"F0";
        when x"3068" => data_out<= x"07";
        when x"3069" => data_out<= x"C6";
        when x"306A" => data_out<= x"0C";
        when x"306B" => data_out<= x"A0";
        when x"306C" => data_out<= x"00";
        when x"306D" => data_out<= x"91";
        when x"306E" => data_out<= x"0C";
        when x"306F" => data_out<= x"60";
        when x"3070" => data_out<= x"C6";
        when x"3071" => data_out<= x"0D";
        when x"3072" => data_out<= x"C6";
        when x"3073" => data_out<= x"0C";
        when x"3074" => data_out<= x"91";
        when x"3075" => data_out<= x"0C";
        when x"3076" => data_out<= x"60";
        when x"3077" => data_out<= x"A9";
        when x"3078" => data_out<= x"00";
        when x"3079" => data_out<= x"A2";
        when x"307A" => data_out<= x"00";
        when x"307B" => data_out<= x"48";
        when x"307C" => data_out<= x"A5";
        when x"307D" => data_out<= x"0C";
        when x"307E" => data_out<= x"38";
        when x"307F" => data_out<= x"E9";
        when x"3080" => data_out<= x"02";
        when x"3081" => data_out<= x"85";
        when x"3082" => data_out<= x"0C";
        when x"3083" => data_out<= x"B0";
        when x"3084" => data_out<= x"02";
        when x"3085" => data_out<= x"C6";
        when x"3086" => data_out<= x"0D";
        when x"3087" => data_out<= x"A0";
        when x"3088" => data_out<= x"01";
        when x"3089" => data_out<= x"8A";
        when x"308A" => data_out<= x"91";
        when x"308B" => data_out<= x"0C";
        when x"308C" => data_out<= x"68";
        when x"308D" => data_out<= x"88";
        when x"308E" => data_out<= x"91";
        when x"308F" => data_out<= x"0C";
        when x"3090" => data_out<= x"60";
        when x"3091" => data_out<= x"A0";
        when x"3092" => data_out<= x"03";
        when x"3093" => data_out<= x"A5";
        when x"3094" => data_out<= x"0C";
        when x"3095" => data_out<= x"38";
        when x"3096" => data_out<= x"E9";
        when x"3097" => data_out<= x"02";
        when x"3098" => data_out<= x"85";
        when x"3099" => data_out<= x"0C";
        when x"309A" => data_out<= x"B0";
        when x"309B" => data_out<= x"02";
        when x"309C" => data_out<= x"C6";
        when x"309D" => data_out<= x"0D";
        when x"309E" => data_out<= x"B1";
        when x"309F" => data_out<= x"0C";
        when x"30A0" => data_out<= x"AA";
        when x"30A1" => data_out<= x"88";
        when x"30A2" => data_out<= x"B1";
        when x"30A3" => data_out<= x"0C";
        when x"30A4" => data_out<= x"A0";
        when x"30A5" => data_out<= x"00";
        when x"30A6" => data_out<= x"91";
        when x"30A7" => data_out<= x"0C";
        when x"30A8" => data_out<= x"C8";
        when x"30A9" => data_out<= x"8A";
        when x"30AA" => data_out<= x"91";
        when x"30AB" => data_out<= x"0C";
        when x"30AC" => data_out<= x"60";
        when x"30AD" => data_out<= x"48";
        when x"30AE" => data_out<= x"84";
        when x"30AF" => data_out<= x"1C";
        when x"30B0" => data_out<= x"A0";
        when x"30B1" => data_out<= x"01";
        when x"30B2" => data_out<= x"B1";
        when x"30B3" => data_out<= x"0C";
        when x"30B4" => data_out<= x"85";
        when x"30B5" => data_out<= x"15";
        when x"30B6" => data_out<= x"88";
        when x"30B7" => data_out<= x"B1";
        when x"30B8" => data_out<= x"0C";
        when x"30B9" => data_out<= x"85";
        when x"30BA" => data_out<= x"14";
        when x"30BB" => data_out<= x"A4";
        when x"30BC" => data_out<= x"1C";
        when x"30BD" => data_out<= x"68";
        when x"30BE" => data_out<= x"91";
        when x"30BF" => data_out<= x"14";
        when x"30C0" => data_out<= x"4C";
        when x"30C1" => data_out<= x"14";
        when x"30C2" => data_out<= x"AF";
        when x"30C3" => data_out<= x"A0";
        when x"30C4" => data_out<= x"00";
        when x"30C5" => data_out<= x"91";
        when x"30C6" => data_out<= x"0C";
        when x"30C7" => data_out<= x"C8";
        when x"30C8" => data_out<= x"48";
        when x"30C9" => data_out<= x"8A";
        when x"30CA" => data_out<= x"91";
        when x"30CB" => data_out<= x"0C";
        when x"30CC" => data_out<= x"68";
        when x"30CD" => data_out<= x"60";
        when x"30CE" => data_out<= x"84";
        when x"30CF" => data_out<= x"1C";
        when x"30D0" => data_out<= x"48";
        when x"30D1" => data_out<= x"A0";
        when x"30D2" => data_out<= x"01";
        when x"30D3" => data_out<= x"B1";
        when x"30D4" => data_out<= x"0C";
        when x"30D5" => data_out<= x"85";
        when x"30D6" => data_out<= x"15";
        when x"30D7" => data_out<= x"88";
        when x"30D8" => data_out<= x"B1";
        when x"30D9" => data_out<= x"0C";
        when x"30DA" => data_out<= x"85";
        when x"30DB" => data_out<= x"14";
        when x"30DC" => data_out<= x"A4";
        when x"30DD" => data_out<= x"1C";
        when x"30DE" => data_out<= x"C8";
        when x"30DF" => data_out<= x"8A";
        when x"30E0" => data_out<= x"91";
        when x"30E1" => data_out<= x"14";
        when x"30E2" => data_out<= x"88";
        when x"30E3" => data_out<= x"68";
        when x"30E4" => data_out<= x"91";
        when x"30E5" => data_out<= x"14";
        when x"30E6" => data_out<= x"4C";
        when x"30E7" => data_out<= x"14";
        when x"30E8" => data_out<= x"AF";
        when x"30E9" => data_out<= x"A0";
        when x"30EA" => data_out<= x"00";
        when x"30EB" => data_out<= x"91";
        when x"30EC" => data_out<= x"0C";
        when x"30ED" => data_out<= x"C8";
        when x"30EE" => data_out<= x"48";
        when x"30EF" => data_out<= x"8A";
        when x"30F0" => data_out<= x"91";
        when x"30F1" => data_out<= x"0C";
        when x"30F2" => data_out<= x"C8";
        when x"30F3" => data_out<= x"A5";
        when x"30F4" => data_out<= x"0E";
        when x"30F5" => data_out<= x"91";
        when x"30F6" => data_out<= x"0C";
        when x"30F7" => data_out<= x"C8";
        when x"30F8" => data_out<= x"A5";
        when x"30F9" => data_out<= x"0F";
        when x"30FA" => data_out<= x"91";
        when x"30FB" => data_out<= x"0C";
        when x"30FC" => data_out<= x"68";
        when x"30FD" => data_out<= x"60";
        when x"30FE" => data_out<= x"A0";
        when x"30FF" => data_out<= x"00";
        when x"3100" => data_out<= x"38";
        when x"3101" => data_out<= x"49";
        when x"3102" => data_out<= x"FF";
        when x"3103" => data_out<= x"71";
        when x"3104" => data_out<= x"0C";
        when x"3105" => data_out<= x"91";
        when x"3106" => data_out<= x"0C";
        when x"3107" => data_out<= x"48";
        when x"3108" => data_out<= x"C8";
        when x"3109" => data_out<= x"8A";
        when x"310A" => data_out<= x"49";
        when x"310B" => data_out<= x"FF";
        when x"310C" => data_out<= x"71";
        when x"310D" => data_out<= x"0C";
        when x"310E" => data_out<= x"91";
        when x"310F" => data_out<= x"0C";
        when x"3110" => data_out<= x"AA";
        when x"3111" => data_out<= x"68";
        when x"3112" => data_out<= x"60";
        when x"3113" => data_out<= x"98";
        when x"3114" => data_out<= x"49";
        when x"3115" => data_out<= x"FF";
        when x"3116" => data_out<= x"38";
        when x"3117" => data_out<= x"65";
        when x"3118" => data_out<= x"0C";
        when x"3119" => data_out<= x"85";
        when x"311A" => data_out<= x"0C";
        when x"311B" => data_out<= x"B0";
        when x"311C" => data_out<= x"02";
        when x"311D" => data_out<= x"C6";
        when x"311E" => data_out<= x"0D";
        when x"311F" => data_out<= x"60";
        when x"3120" => data_out<= x"A2";
        when x"3121" => data_out<= x"00";
        when x"3122" => data_out<= x"85";
        when x"3123" => data_out<= x"1A";
        when x"3124" => data_out<= x"86";
        when x"3125" => data_out<= x"1B";
        when x"3126" => data_out<= x"20";
        when x"3127" => data_out<= x"53";
        when x"3128" => data_out<= x"B0";
        when x"3129" => data_out<= x"20";
        when x"312A" => data_out<= x"31";
        when x"312B" => data_out<= x"B1";
        when x"312C" => data_out<= x"A5";
        when x"312D" => data_out<= x"14";
        when x"312E" => data_out<= x"A6";
        when x"312F" => data_out<= x"15";
        when x"3130" => data_out<= x"60";
        when x"3131" => data_out<= x"A9";
        when x"3132" => data_out<= x"00";
        when x"3133" => data_out<= x"85";
        when x"3134" => data_out<= x"0F";
        when x"3135" => data_out<= x"A0";
        when x"3136" => data_out<= x"10";
        when x"3137" => data_out<= x"A6";
        when x"3138" => data_out<= x"1B";
        when x"3139" => data_out<= x"F0";
        when x"313A" => data_out<= x"1F";
        when x"313B" => data_out<= x"06";
        when x"313C" => data_out<= x"14";
        when x"313D" => data_out<= x"26";
        when x"313E" => data_out<= x"15";
        when x"313F" => data_out<= x"2A";
        when x"3140" => data_out<= x"26";
        when x"3141" => data_out<= x"0F";
        when x"3142" => data_out<= x"AA";
        when x"3143" => data_out<= x"C5";
        when x"3144" => data_out<= x"1A";
        when x"3145" => data_out<= x"A5";
        when x"3146" => data_out<= x"0F";
        when x"3147" => data_out<= x"E5";
        when x"3148" => data_out<= x"1B";
        when x"3149" => data_out<= x"90";
        when x"314A" => data_out<= x"08";
        when x"314B" => data_out<= x"85";
        when x"314C" => data_out<= x"0F";
        when x"314D" => data_out<= x"8A";
        when x"314E" => data_out<= x"E5";
        when x"314F" => data_out<= x"1A";
        when x"3150" => data_out<= x"AA";
        when x"3151" => data_out<= x"E6";
        when x"3152" => data_out<= x"14";
        when x"3153" => data_out<= x"8A";
        when x"3154" => data_out<= x"88";
        when x"3155" => data_out<= x"D0";
        when x"3156" => data_out<= x"E4";
        when x"3157" => data_out<= x"85";
        when x"3158" => data_out<= x"0E";
        when x"3159" => data_out<= x"60";
        when x"315A" => data_out<= x"06";
        when x"315B" => data_out<= x"14";
        when x"315C" => data_out<= x"26";
        when x"315D" => data_out<= x"15";
        when x"315E" => data_out<= x"2A";
        when x"315F" => data_out<= x"B0";
        when x"3160" => data_out<= x"04";
        when x"3161" => data_out<= x"C5";
        when x"3162" => data_out<= x"1A";
        when x"3163" => data_out<= x"90";
        when x"3164" => data_out<= x"04";
        when x"3165" => data_out<= x"E5";
        when x"3166" => data_out<= x"1A";
        when x"3167" => data_out<= x"E6";
        when x"3168" => data_out<= x"14";
        when x"3169" => data_out<= x"88";
        when x"316A" => data_out<= x"D0";
        when x"316B" => data_out<= x"EE";
        when x"316C" => data_out<= x"85";
        when x"316D" => data_out<= x"0E";
        when x"316E" => data_out<= x"60";
        when x"316F" => data_out<= x"A2";
        when x"3170" => data_out<= x"00";
        when x"3171" => data_out<= x"85";
        when x"3172" => data_out<= x"1A";
        when x"3173" => data_out<= x"86";
        when x"3174" => data_out<= x"1B";
        when x"3175" => data_out<= x"20";
        when x"3176" => data_out<= x"53";
        when x"3177" => data_out<= x"B0";
        when x"3178" => data_out<= x"20";
        when x"3179" => data_out<= x"31";
        when x"317A" => data_out<= x"B1";
        when x"317B" => data_out<= x"A5";
        when x"317C" => data_out<= x"0E";
        when x"317D" => data_out<= x"A6";
        when x"317E" => data_out<= x"0F";
        when x"317F" => data_out<= x"60";
        when x"3180" => data_out<= x"23";
        when x"3181" => data_out<= x"23";
        when x"3182" => data_out<= x"23";
        when x"3183" => data_out<= x"23";
        when x"3184" => data_out<= x"23";
        when x"3185" => data_out<= x"20";
        when x"3186" => data_out<= x"36";
        when x"3187" => data_out<= x"35";
        when x"3188" => data_out<= x"30";
        when x"3189" => data_out<= x"32";
        when x"318A" => data_out<= x"20";
        when x"318B" => data_out<= x"53";
        when x"318C" => data_out<= x"59";
        when x"318D" => data_out<= x"53";
        when x"318E" => data_out<= x"54";
        when x"318F" => data_out<= x"45";
        when x"3190" => data_out<= x"4D";
        when x"3191" => data_out<= x"20";
        when x"3192" => data_out<= x"52";
        when x"3193" => data_out<= x"45";
        when x"3194" => data_out<= x"41";
        when x"3195" => data_out<= x"44";
        when x"3196" => data_out<= x"59";
        when x"3197" => data_out<= x"20";
        when x"3198" => data_out<= x"23";
        when x"3199" => data_out<= x"23";
        when x"319A" => data_out<= x"23";
        when x"319B" => data_out<= x"23";
        when x"319C" => data_out<= x"23";
        when x"319D" => data_out<= x"0D";
        when x"319E" => data_out<= x"0A";
        when x"319F" => data_out<= x"00";
        when x"31A0" => data_out<= x"52";
        when x"31A1" => data_out<= x"65";
        when x"31A2" => data_out<= x"69";
        when x"31A3" => data_out<= x"6E";
        when x"31A4" => data_out<= x"69";
        when x"31A5" => data_out<= x"63";
        when x"31A6" => data_out<= x"69";
        when x"31A7" => data_out<= x"61";
        when x"31A8" => data_out<= x"6E";
        when x"31A9" => data_out<= x"64";
        when x"31AA" => data_out<= x"6F";
        when x"31AB" => data_out<= x"20";
        when x"31AC" => data_out<= x"6D";
        when x"31AD" => data_out<= x"6F";
        when x"31AE" => data_out<= x"6E";
        when x"31AF" => data_out<= x"69";
        when x"31B0" => data_out<= x"74";
        when x"31B1" => data_out<= x"6F";
        when x"31B2" => data_out<= x"72";
        when x"31B3" => data_out<= x"2E";
        when x"31B4" => data_out<= x"2E";
        when x"31B5" => data_out<= x"2E";
        when x"31B6" => data_out<= x"0D";
        when x"31B7" => data_out<= x"0A";
        when x"31B8" => data_out<= x"00";
        when x"31B9" => data_out<= x"49";
        when x"31BA" => data_out<= x"6E";
        when x"31BB" => data_out<= x"69";
        when x"31BC" => data_out<= x"63";
        when x"31BD" => data_out<= x"69";
        when x"31BE" => data_out<= x"61";
        when x"31BF" => data_out<= x"6E";
        when x"31C0" => data_out<= x"64";
        when x"31C1" => data_out<= x"6F";
        when x"31C2" => data_out<= x"20";
        when x"31C3" => data_out<= x"4D";
        when x"31C4" => data_out<= x"6F";
        when x"31C5" => data_out<= x"6E";
        when x"31C6" => data_out<= x"69";
        when x"31C7" => data_out<= x"74";
        when x"31C8" => data_out<= x"6F";
        when x"31C9" => data_out<= x"72";
        when x"31CA" => data_out<= x"2E";
        when x"31CB" => data_out<= x"2E";
        when x"31CC" => data_out<= x"2E";
        when x"31CD" => data_out<= x"0D";
        when x"31CE" => data_out<= x"0A";
        when x"31CF" => data_out<= x"00";
        when x"31D0" => data_out<= x"30";
        when x"31D1" => data_out<= x"31";
        when x"31D2" => data_out<= x"32";
        when x"31D3" => data_out<= x"33";
        when x"31D4" => data_out<= x"34";
        when x"31D5" => data_out<= x"35";
        when x"31D6" => data_out<= x"36";
        when x"31D7" => data_out<= x"37";
        when x"31D8" => data_out<= x"38";
        when x"31D9" => data_out<= x"39";
        when x"31DA" => data_out<= x"41";
        when x"31DB" => data_out<= x"42";
        when x"31DC" => data_out<= x"43";
        when x"31DD" => data_out<= x"44";
        when x"31DE" => data_out<= x"45";
        when x"31DF" => data_out<= x"46";
        when x"31E0" => data_out<= x"00";
        when x"31E1" => data_out<= x"43";
        when x"31E2" => data_out<= x"6D";
        when x"31E3" => data_out<= x"64";
        when x"31E4" => data_out<= x"73";
        when x"31E5" => data_out<= x"20";
        when x"31E6" => data_out<= x"53";
        when x"31E7" => data_out<= x"44";
        when x"31E8" => data_out<= x"3A";
        when x"31E9" => data_out<= x"20";
        when x"31EA" => data_out<= x"53";
        when x"31EB" => data_out<= x"44";
        when x"31EC" => data_out<= x"2C";
        when x"31ED" => data_out<= x"4C";
        when x"31EE" => data_out<= x"53";
        when x"31EF" => data_out<= x"2C";
        when x"31F0" => data_out<= x"53";
        when x"31F1" => data_out<= x"41";
        when x"31F2" => data_out<= x"56";
        when x"31F3" => data_out<= x"45";
        when x"31F4" => data_out<= x"2C";
        when x"31F5" => data_out<= x"4C";
        when x"31F6" => data_out<= x"4F";
        when x"31F7" => data_out<= x"41";
        when x"31F8" => data_out<= x"44";
        when x"31F9" => data_out<= x"2C";
        when x"31FA" => data_out<= x"44";
        when x"31FB" => data_out<= x"45";
        when x"31FC" => data_out<= x"4C";
        when x"31FD" => data_out<= x"2C";
        when x"31FE" => data_out<= x"43";
        when x"31FF" => data_out<= x"41";
        when x"3200" => data_out<= x"54";
        when x"3201" => data_out<= x"2C";
        when x"3202" => data_out<= x"53";
        when x"3203" => data_out<= x"44";
        when x"3204" => data_out<= x"46";
        when x"3205" => data_out<= x"4F";
        when x"3206" => data_out<= x"52";
        when x"3207" => data_out<= x"4D";
        when x"3208" => data_out<= x"41";
        when x"3209" => data_out<= x"54";
        when x"320A" => data_out<= x"0D";
        when x"320B" => data_out<= x"0A";
        when x"320C" => data_out<= x"00";
        when x"320D" => data_out<= x"4D";
        when x"320E" => data_out<= x"75";
        when x"320F" => data_out<= x"65";
        when x"3210" => data_out<= x"73";
        when x"3211" => data_out<= x"74";
        when x"3212" => data_out<= x"72";
        when x"3213" => data_out<= x"61";
        when x"3214" => data_out<= x"20";
        when x"3215" => data_out<= x"72";
        when x"3216" => data_out<= x"61";
        when x"3217" => data_out<= x"6E";
        when x"3218" => data_out<= x"67";
        when x"3219" => data_out<= x"6F";
        when x"321A" => data_out<= x"73";
        when x"321B" => data_out<= x"3A";
        when x"321C" => data_out<= x"20";
        when x"321D" => data_out<= x"5A";
        when x"321E" => data_out<= x"50";
        when x"321F" => data_out<= x"2C";
        when x"3220" => data_out<= x"53";
        when x"3221" => data_out<= x"74";
        when x"3222" => data_out<= x"61";
        when x"3223" => data_out<= x"63";
        when x"3224" => data_out<= x"6B";
        when x"3225" => data_out<= x"2C";
        when x"3226" => data_out<= x"52";
        when x"3227" => data_out<= x"41";
        when x"3228" => data_out<= x"4D";
        when x"3229" => data_out<= x"2C";
        when x"322A" => data_out<= x"49";
        when x"322B" => data_out<= x"2F";
        when x"322C" => data_out<= x"4F";
        when x"322D" => data_out<= x"2C";
        when x"322E" => data_out<= x"52";
        when x"322F" => data_out<= x"4F";
        when x"3230" => data_out<= x"4D";
        when x"3231" => data_out<= x"0D";
        when x"3232" => data_out<= x"0A";
        when x"3233" => data_out<= x"00";
        when x"3234" => data_out<= x"45";
        when x"3235" => data_out<= x"73";
        when x"3236" => data_out<= x"63";
        when x"3237" => data_out<= x"72";
        when x"3238" => data_out<= x"69";
        when x"3239" => data_out<= x"62";
        when x"323A" => data_out<= x"65";
        when x"323B" => data_out<= x"20";
        when x"323C" => data_out<= x"48";
        when x"323D" => data_out<= x"20";
        when x"323E" => data_out<= x"70";
        when x"323F" => data_out<= x"61";
        when x"3240" => data_out<= x"72";
        when x"3241" => data_out<= x"61";
        when x"3242" => data_out<= x"20";
        when x"3243" => data_out<= x"61";
        when x"3244" => data_out<= x"79";
        when x"3245" => data_out<= x"75";
        when x"3246" => data_out<= x"64";
        when x"3247" => data_out<= x"61";
        when x"3248" => data_out<= x"2C";
        when x"3249" => data_out<= x"20";
        when x"324A" => data_out<= x"53";
        when x"324B" => data_out<= x"44";
        when x"324C" => data_out<= x"20";
        when x"324D" => data_out<= x"70";
        when x"324E" => data_out<= x"61";
        when x"324F" => data_out<= x"72";
        when x"3250" => data_out<= x"61";
        when x"3251" => data_out<= x"20";
        when x"3252" => data_out<= x"53";
        when x"3253" => data_out<= x"44";
        when x"3254" => data_out<= x"20";
        when x"3255" => data_out<= x"43";
        when x"3256" => data_out<= x"61";
        when x"3257" => data_out<= x"72";
        when x"3258" => data_out<= x"64";
        when x"3259" => data_out<= x"00";
        when x"325A" => data_out<= x"56";
        when x"325B" => data_out<= x"61";
        when x"325C" => data_out<= x"6C";
        when x"325D" => data_out<= x"6F";
        when x"325E" => data_out<= x"72";
        when x"325F" => data_out<= x"65";
        when x"3260" => data_out<= x"73";
        when x"3261" => data_out<= x"20";
        when x"3262" => data_out<= x"48";
        when x"3263" => data_out<= x"45";
        when x"3264" => data_out<= x"58";
        when x"3265" => data_out<= x"2E";
        when x"3266" => data_out<= x"20";
        when x"3267" => data_out<= x"48";
        when x"3268" => data_out<= x"20";
        when x"3269" => data_out<= x"63";
        when x"326A" => data_out<= x"6D";
        when x"326B" => data_out<= x"64";
        when x"326C" => data_out<= x"3D";
        when x"326D" => data_out<= x"61";
        when x"326E" => data_out<= x"79";
        when x"326F" => data_out<= x"75";
        when x"3270" => data_out<= x"64";
        when x"3271" => data_out<= x"61";
        when x"3272" => data_out<= x"20";
        when x"3273" => data_out<= x"64";
        when x"3274" => data_out<= x"65";
        when x"3275" => data_out<= x"74";
        when x"3276" => data_out<= x"61";
        when x"3277" => data_out<= x"6C";
        when x"3278" => data_out<= x"6C";
        when x"3279" => data_out<= x"61";
        when x"327A" => data_out<= x"64";
        when x"327B" => data_out<= x"61";
        when x"327C" => data_out<= x"0D";
        when x"327D" => data_out<= x"0A";
        when x"327E" => data_out<= x"00";
        when x"327F" => data_out<= x"45";
        when x"3280" => data_out<= x"6A";
        when x"3281" => data_out<= x"3A";
        when x"3282" => data_out<= x"20";
        when x"3283" => data_out<= x"4C";
        when x"3284" => data_out<= x"4F";
        when x"3285" => data_out<= x"41";
        when x"3286" => data_out<= x"44";
        when x"3287" => data_out<= x"20";
        when x"3288" => data_out<= x"50";
        when x"3289" => data_out<= x"52";
        when x"328A" => data_out<= x"4F";
        when x"328B" => data_out<= x"47";
        when x"328C" => data_out<= x"2E";
        when x"328D" => data_out<= x"42";
        when x"328E" => data_out<= x"49";
        when x"328F" => data_out<= x"4E";
        when x"3290" => data_out<= x"2C";
        when x"3291" => data_out<= x"20";
        when x"3292" => data_out<= x"4C";
        when x"3293" => data_out<= x"4F";
        when x"3294" => data_out<= x"41";
        when x"3295" => data_out<= x"44";
        when x"3296" => data_out<= x"20";
        when x"3297" => data_out<= x"50";
        when x"3298" => data_out<= x"2E";
        when x"3299" => data_out<= x"42";
        when x"329A" => data_out<= x"49";
        when x"329B" => data_out<= x"4E";
        when x"329C" => data_out<= x"20";
        when x"329D" => data_out<= x"31";
        when x"329E" => data_out<= x"30";
        when x"329F" => data_out<= x"30";
        when x"32A0" => data_out<= x"30";
        when x"32A1" => data_out<= x"0D";
        when x"32A2" => data_out<= x"0A";
        when x"32A3" => data_out<= x"00";
        when x"32A4" => data_out<= x"45";
        when x"32A5" => data_out<= x"6A";
        when x"32A6" => data_out<= x"3A";
        when x"32A7" => data_out<= x"20";
        when x"32A8" => data_out<= x"4C";
        when x"32A9" => data_out<= x"20";
        when x"32AA" => data_out<= x"30";
        when x"32AB" => data_out<= x"32";
        when x"32AC" => data_out<= x"30";
        when x"32AD" => data_out<= x"30";
        when x"32AE" => data_out<= x"20";
        when x"32AF" => data_out<= x"2D";
        when x"32B0" => data_out<= x"3E";
        when x"32B1" => data_out<= x"20";
        when x"32B2" => data_out<= x"41";
        when x"32B3" => data_out<= x"39";
        when x"32B4" => data_out<= x"20";
        when x"32B5" => data_out<= x"30";
        when x"32B6" => data_out<= x"31";
        when x"32B7" => data_out<= x"20";
        when x"32B8" => data_out<= x"38";
        when x"32B9" => data_out<= x"44";
        when x"32BA" => data_out<= x"20";
        when x"32BB" => data_out<= x"30";
        when x"32BC" => data_out<= x"31";
        when x"32BD" => data_out<= x"20";
        when x"32BE" => data_out<= x"43";
        when x"32BF" => data_out<= x"30";
        when x"32C0" => data_out<= x"20";
        when x"32C1" => data_out<= x"36";
        when x"32C2" => data_out<= x"30";
        when x"32C3" => data_out<= x"20";
        when x"32C4" => data_out<= x"2E";
        when x"32C5" => data_out<= x"0D";
        when x"32C6" => data_out<= x"0A";
        when x"32C7" => data_out<= x"00";
        when x"32C8" => data_out<= x"53";
        when x"32C9" => data_out<= x"44";
        when x"32CA" => data_out<= x"2F";
        when x"32CB" => data_out<= x"4C";
        when x"32CC" => data_out<= x"53";
        when x"32CD" => data_out<= x"2F";
        when x"32CE" => data_out<= x"53";
        when x"32CF" => data_out<= x"44";
        when x"32D0" => data_out<= x"46";
        when x"32D1" => data_out<= x"4F";
        when x"32D2" => data_out<= x"52";
        when x"32D3" => data_out<= x"4D";
        when x"32D4" => data_out<= x"41";
        when x"32D5" => data_out<= x"54";
        when x"32D6" => data_out<= x"20";
        when x"32D7" => data_out<= x"53";
        when x"32D8" => data_out<= x"41";
        when x"32D9" => data_out<= x"56";
        when x"32DA" => data_out<= x"45";
        when x"32DB" => data_out<= x"2F";
        when x"32DC" => data_out<= x"4C";
        when x"32DD" => data_out<= x"4F";
        when x"32DE" => data_out<= x"41";
        when x"32DF" => data_out<= x"44";
        when x"32E0" => data_out<= x"2F";
        when x"32E1" => data_out<= x"44";
        when x"32E2" => data_out<= x"45";
        when x"32E3" => data_out<= x"4C";
        when x"32E4" => data_out<= x"2F";
        when x"32E5" => data_out<= x"43";
        when x"32E6" => data_out<= x"41";
        when x"32E7" => data_out<= x"54";
        when x"32E8" => data_out<= x"0D";
        when x"32E9" => data_out<= x"0A";
        when x"32EA" => data_out<= x"00";
        when x"32EB" => data_out<= x"4C";
        when x"32EC" => data_out<= x"20";
        when x"32ED" => data_out<= x"61";
        when x"32EE" => data_out<= x"64";
        when x"32EF" => data_out<= x"64";
        when x"32F0" => data_out<= x"72";
        when x"32F1" => data_out<= x"20";
        when x"32F2" => data_out<= x"2D";
        when x"32F3" => data_out<= x"20";
        when x"32F4" => data_out<= x"43";
        when x"32F5" => data_out<= x"61";
        when x"32F6" => data_out<= x"72";
        when x"32F7" => data_out<= x"67";
        when x"32F8" => data_out<= x"61";
        when x"32F9" => data_out<= x"72";
        when x"32FA" => data_out<= x"20";
        when x"32FB" => data_out<= x"68";
        when x"32FC" => data_out<= x"65";
        when x"32FD" => data_out<= x"78";
        when x"32FE" => data_out<= x"20";
        when x"32FF" => data_out<= x"69";
        when x"3300" => data_out<= x"6E";
        when x"3301" => data_out<= x"74";
        when x"3302" => data_out<= x"65";
        when x"3303" => data_out<= x"72";
        when x"3304" => data_out<= x"61";
        when x"3305" => data_out<= x"63";
        when x"3306" => data_out<= x"74";
        when x"3307" => data_out<= x"69";
        when x"3308" => data_out<= x"76";
        when x"3309" => data_out<= x"6F";
        when x"330A" => data_out<= x"0D";
        when x"330B" => data_out<= x"0A";
        when x"330C" => data_out<= x"00";
        when x"330D" => data_out<= x"58";
        when x"330E" => data_out<= x"52";
        when x"330F" => data_out<= x"45";
        when x"3310" => data_out<= x"43";
        when x"3311" => data_out<= x"56";
        when x"3312" => data_out<= x"20";
        when x"3313" => data_out<= x"5B";
        when x"3314" => data_out<= x"61";
        when x"3315" => data_out<= x"64";
        when x"3316" => data_out<= x"64";
        when x"3317" => data_out<= x"72";
        when x"3318" => data_out<= x"5D";
        when x"3319" => data_out<= x"20";
        when x"331A" => data_out<= x"58";
        when x"331B" => data_out<= x"4D";
        when x"331C" => data_out<= x"4F";
        when x"331D" => data_out<= x"44";
        when x"331E" => data_out<= x"45";
        when x"331F" => data_out<= x"4D";
        when x"3320" => data_out<= x"20";
        when x"3321" => data_out<= x"28";
        when x"3322" => data_out<= x"64";
        when x"3323" => data_out<= x"65";
        when x"3324" => data_out<= x"66";
        when x"3325" => data_out<= x"20";
        when x"3326" => data_out<= x"24";
        when x"3327" => data_out<= x"30";
        when x"3328" => data_out<= x"38";
        when x"3329" => data_out<= x"30";
        when x"332A" => data_out<= x"30";
        when x"332B" => data_out<= x"29";
        when x"332C" => data_out<= x"0D";
        when x"332D" => data_out<= x"0A";
        when x"332E" => data_out<= x"00";
        when x"332F" => data_out<= x"45";
        when x"3330" => data_out<= x"6A";
        when x"3331" => data_out<= x"3A";
        when x"3332" => data_out<= x"20";
        when x"3333" => data_out<= x"46";
        when x"3334" => data_out<= x"20";
        when x"3335" => data_out<= x"30";
        when x"3336" => data_out<= x"32";
        when x"3337" => data_out<= x"30";
        when x"3338" => data_out<= x"30";
        when x"3339" => data_out<= x"20";
        when x"333A" => data_out<= x"31";
        when x"333B" => data_out<= x"30";
        when x"333C" => data_out<= x"30";
        when x"333D" => data_out<= x"20";
        when x"333E" => data_out<= x"30";
        when x"333F" => data_out<= x"30";
        when x"3340" => data_out<= x"2C";
        when x"3341" => data_out<= x"20";
        when x"3342" => data_out<= x"46";
        when x"3343" => data_out<= x"20";
        when x"3344" => data_out<= x"30";
        when x"3345" => data_out<= x"32";
        when x"3346" => data_out<= x"30";
        when x"3347" => data_out<= x"30";
        when x"3348" => data_out<= x"20";
        when x"3349" => data_out<= x"31";
        when x"334A" => data_out<= x"30";
        when x"334B" => data_out<= x"20";
        when x"334C" => data_out<= x"45";
        when x"334D" => data_out<= x"41";
        when x"334E" => data_out<= x"0D";
        when x"334F" => data_out<= x"0A";
        when x"3350" => data_out<= x"00";
        when x"3351" => data_out<= x"6C";
        when x"3352" => data_out<= x"65";
        when x"3353" => data_out<= x"6E";
        when x"3354" => data_out<= x"20";
        when x"3355" => data_out<= x"64";
        when x"3356" => data_out<= x"65";
        when x"3357" => data_out<= x"66";
        when x"3358" => data_out<= x"61";
        when x"3359" => data_out<= x"75";
        when x"335A" => data_out<= x"6C";
        when x"335B" => data_out<= x"74";
        when x"335C" => data_out<= x"3D";
        when x"335D" => data_out<= x"36";
        when x"335E" => data_out<= x"34";
        when x"335F" => data_out<= x"2E";
        when x"3360" => data_out<= x"20";
        when x"3361" => data_out<= x"45";
        when x"3362" => data_out<= x"6A";
        when x"3363" => data_out<= x"3A";
        when x"3364" => data_out<= x"20";
        when x"3365" => data_out<= x"44";
        when x"3366" => data_out<= x"20";
        when x"3367" => data_out<= x"30";
        when x"3368" => data_out<= x"32";
        when x"3369" => data_out<= x"30";
        when x"336A" => data_out<= x"30";
        when x"336B" => data_out<= x"20";
        when x"336C" => data_out<= x"31";
        when x"336D" => data_out<= x"30";
        when x"336E" => data_out<= x"30";
        when x"336F" => data_out<= x"0D";
        when x"3370" => data_out<= x"0A";
        when x"3371" => data_out<= x"00";
        when x"3372" => data_out<= x"45";
        when x"3373" => data_out<= x"6A";
        when x"3374" => data_out<= x"65";
        when x"3375" => data_out<= x"63";
        when x"3376" => data_out<= x"75";
        when x"3377" => data_out<= x"74";
        when x"3378" => data_out<= x"61";
        when x"3379" => data_out<= x"72";
        when x"337A" => data_out<= x"20";
        when x"337B" => data_out<= x"61";
        when x"337C" => data_out<= x"6E";
        when x"337D" => data_out<= x"74";
        when x"337E" => data_out<= x"65";
        when x"337F" => data_out<= x"73";
        when x"3380" => data_out<= x"20";
        when x"3381" => data_out<= x"64";
        when x"3382" => data_out<= x"65";
        when x"3383" => data_out<= x"20";
        when x"3384" => data_out<= x"6F";
        when x"3385" => data_out<= x"74";
        when x"3386" => data_out<= x"72";
        when x"3387" => data_out<= x"6F";
        when x"3388" => data_out<= x"73";
        when x"3389" => data_out<= x"20";
        when x"338A" => data_out<= x"63";
        when x"338B" => data_out<= x"6D";
        when x"338C" => data_out<= x"64";
        when x"338D" => data_out<= x"20";
        when x"338E" => data_out<= x"53";
        when x"338F" => data_out<= x"44";
        when x"3390" => data_out<= x"0D";
        when x"3391" => data_out<= x"0A";
        when x"3392" => data_out<= x"00";
        when x"3393" => data_out<= x"3D";
        when x"3394" => data_out<= x"3D";
        when x"3395" => data_out<= x"3D";
        when x"3396" => data_out<= x"3D";
        when x"3397" => data_out<= x"3D";
        when x"3398" => data_out<= x"3D";
        when x"3399" => data_out<= x"3D";
        when x"339A" => data_out<= x"3D";
        when x"339B" => data_out<= x"3D";
        when x"339C" => data_out<= x"3D";
        when x"339D" => data_out<= x"3D";
        when x"339E" => data_out<= x"3D";
        when x"339F" => data_out<= x"3D";
        when x"33A0" => data_out<= x"3D";
        when x"33A1" => data_out<= x"3D";
        when x"33A2" => data_out<= x"3D";
        when x"33A3" => data_out<= x"3D";
        when x"33A4" => data_out<= x"3D";
        when x"33A5" => data_out<= x"3D";
        when x"33A6" => data_out<= x"3D";
        when x"33A7" => data_out<= x"3D";
        when x"33A8" => data_out<= x"3D";
        when x"33A9" => data_out<= x"3D";
        when x"33AA" => data_out<= x"3D";
        when x"33AB" => data_out<= x"3D";
        when x"33AC" => data_out<= x"3D";
        when x"33AD" => data_out<= x"3D";
        when x"33AE" => data_out<= x"3D";
        when x"33AF" => data_out<= x"3D";
        when x"33B0" => data_out<= x"3D";
        when x"33B1" => data_out<= x"3D";
        when x"33B2" => data_out<= x"3D";
        when x"33B3" => data_out<= x"00";
        when x"33B4" => data_out<= x"52";
        when x"33B5" => data_out<= x"20";
        when x"33B6" => data_out<= x"5B";
        when x"33B7" => data_out<= x"61";
        when x"33B8" => data_out<= x"64";
        when x"33B9" => data_out<= x"64";
        when x"33BA" => data_out<= x"72";
        when x"33BB" => data_out<= x"5D";
        when x"33BC" => data_out<= x"20";
        when x"33BD" => data_out<= x"2D";
        when x"33BE" => data_out<= x"20";
        when x"33BF" => data_out<= x"52";
        when x"33C0" => data_out<= x"75";
        when x"33C1" => data_out<= x"6E";
        when x"33C2" => data_out<= x"2F";
        when x"33C3" => data_out<= x"65";
        when x"33C4" => data_out<= x"6A";
        when x"33C5" => data_out<= x"65";
        when x"33C6" => data_out<= x"63";
        when x"33C7" => data_out<= x"75";
        when x"33C8" => data_out<= x"74";
        when x"33C9" => data_out<= x"61";
        when x"33CA" => data_out<= x"72";
        when x"33CB" => data_out<= x"20";
        when x"33CC" => data_out<= x"63";
        when x"33CD" => data_out<= x"6F";
        when x"33CE" => data_out<= x"64";
        when x"33CF" => data_out<= x"69";
        when x"33D0" => data_out<= x"67";
        when x"33D1" => data_out<= x"6F";
        when x"33D2" => data_out<= x"0D";
        when x"33D3" => data_out<= x"0A";
        when x"33D4" => data_out<= x"00";
        when x"33D5" => data_out<= x"44";
        when x"33D6" => data_out<= x"20";
        when x"33D7" => data_out<= x"61";
        when x"33D8" => data_out<= x"64";
        when x"33D9" => data_out<= x"64";
        when x"33DA" => data_out<= x"72";
        when x"33DB" => data_out<= x"20";
        when x"33DC" => data_out<= x"5B";
        when x"33DD" => data_out<= x"6C";
        when x"33DE" => data_out<= x"65";
        when x"33DF" => data_out<= x"6E";
        when x"33E0" => data_out<= x"5D";
        when x"33E1" => data_out<= x"20";
        when x"33E2" => data_out<= x"2D";
        when x"33E3" => data_out<= x"20";
        when x"33E4" => data_out<= x"44";
        when x"33E5" => data_out<= x"75";
        when x"33E6" => data_out<= x"6D";
        when x"33E7" => data_out<= x"70";
        when x"33E8" => data_out<= x"20";
        when x"33E9" => data_out<= x"68";
        when x"33EA" => data_out<= x"65";
        when x"33EB" => data_out<= x"78";
        when x"33EC" => data_out<= x"2B";
        when x"33ED" => data_out<= x"41";
        when x"33EE" => data_out<= x"53";
        when x"33EF" => data_out<= x"43";
        when x"33F0" => data_out<= x"49";
        when x"33F1" => data_out<= x"49";
        when x"33F2" => data_out<= x"0D";
        when x"33F3" => data_out<= x"0A";
        when x"33F4" => data_out<= x"00";
        when x"33F5" => data_out<= x"52";
        when x"33F6" => data_out<= x"4F";
        when x"33F7" => data_out<= x"4D";
        when x"33F8" => data_out<= x"3A";
        when x"33F9" => data_out<= x"20";
        when x"33FA" => data_out<= x"20";
        when x"33FB" => data_out<= x"20";
        when x"33FC" => data_out<= x"20";
        when x"33FD" => data_out<= x"20";
        when x"33FE" => data_out<= x"20";
        when x"33FF" => data_out<= x"20";
        when x"3400" => data_out<= x"20";
        when x"3401" => data_out<= x"24";
        when x"3402" => data_out<= x"38";
        when x"3403" => data_out<= x"30";
        when x"3404" => data_out<= x"30";
        when x"3405" => data_out<= x"30";
        when x"3406" => data_out<= x"2D";
        when x"3407" => data_out<= x"24";
        when x"3408" => data_out<= x"42";
        when x"3409" => data_out<= x"46";
        when x"340A" => data_out<= x"46";
        when x"340B" => data_out<= x"46";
        when x"340C" => data_out<= x"20";
        when x"340D" => data_out<= x"28";
        when x"340E" => data_out<= x"31";
        when x"340F" => data_out<= x"36";
        when x"3410" => data_out<= x"20";
        when x"3411" => data_out<= x"4B";
        when x"3412" => data_out<= x"42";
        when x"3413" => data_out<= x"29";
        when x"3414" => data_out<= x"00";
        when x"3415" => data_out<= x"46";
        when x"3416" => data_out<= x"20";
        when x"3417" => data_out<= x"61";
        when x"3418" => data_out<= x"64";
        when x"3419" => data_out<= x"64";
        when x"341A" => data_out<= x"72";
        when x"341B" => data_out<= x"20";
        when x"341C" => data_out<= x"6C";
        when x"341D" => data_out<= x"65";
        when x"341E" => data_out<= x"6E";
        when x"341F" => data_out<= x"20";
        when x"3420" => data_out<= x"76";
        when x"3421" => data_out<= x"61";
        when x"3422" => data_out<= x"6C";
        when x"3423" => data_out<= x"20";
        when x"3424" => data_out<= x"2D";
        when x"3425" => data_out<= x"20";
        when x"3426" => data_out<= x"46";
        when x"3427" => data_out<= x"69";
        when x"3428" => data_out<= x"6C";
        when x"3429" => data_out<= x"6C";
        when x"342A" => data_out<= x"20";
        when x"342B" => data_out<= x"6D";
        when x"342C" => data_out<= x"65";
        when x"342D" => data_out<= x"6D";
        when x"342E" => data_out<= x"6F";
        when x"342F" => data_out<= x"72";
        when x"3430" => data_out<= x"69";
        when x"3431" => data_out<= x"61";
        when x"3432" => data_out<= x"0D";
        when x"3433" => data_out<= x"0A";
        when x"3434" => data_out<= x"00";
        when x"3435" => data_out<= x"58";
        when x"3436" => data_out<= x"52";
        when x"3437" => data_out<= x"45";
        when x"3438" => data_out<= x"43";
        when x"3439" => data_out<= x"56";
        when x"343A" => data_out<= x"20";
        when x"343B" => data_out<= x"5B";
        when x"343C" => data_out<= x"61";
        when x"343D" => data_out<= x"64";
        when x"343E" => data_out<= x"64";
        when x"343F" => data_out<= x"72";
        when x"3440" => data_out<= x"5D";
        when x"3441" => data_out<= x"20";
        when x"3442" => data_out<= x"2D";
        when x"3443" => data_out<= x"20";
        when x"3444" => data_out<= x"52";
        when x"3445" => data_out<= x"65";
        when x"3446" => data_out<= x"63";
        when x"3447" => data_out<= x"69";
        when x"3448" => data_out<= x"62";
        when x"3449" => data_out<= x"69";
        when x"344A" => data_out<= x"72";
        when x"344B" => data_out<= x"20";
        when x"344C" => data_out<= x"58";
        when x"344D" => data_out<= x"4D";
        when x"344E" => data_out<= x"4F";
        when x"344F" => data_out<= x"44";
        when x"3450" => data_out<= x"45";
        when x"3451" => data_out<= x"4D";
        when x"3452" => data_out<= x"0D";
        when x"3453" => data_out<= x"0A";
        when x"3454" => data_out<= x"00";
        when x"3455" => data_out<= x"4C";
        when x"3456" => data_out<= x"20";
        when x"3457" => data_out<= x"61";
        when x"3458" => data_out<= x"64";
        when x"3459" => data_out<= x"64";
        when x"345A" => data_out<= x"72";
        when x"345B" => data_out<= x"20";
        when x"345C" => data_out<= x"20";
        when x"345D" => data_out<= x"20";
        when x"345E" => data_out<= x"20";
        when x"345F" => data_out<= x"20";
        when x"3460" => data_out<= x"43";
        when x"3461" => data_out<= x"61";
        when x"3462" => data_out<= x"72";
        when x"3463" => data_out<= x"67";
        when x"3464" => data_out<= x"61";
        when x"3465" => data_out<= x"72";
        when x"3466" => data_out<= x"20";
        when x"3467" => data_out<= x"68";
        when x"3468" => data_out<= x"65";
        when x"3469" => data_out<= x"78";
        when x"346A" => data_out<= x"28";
        when x"346B" => data_out<= x"2E";
        when x"346C" => data_out<= x"3D";
        when x"346D" => data_out<= x"66";
        when x"346E" => data_out<= x"69";
        when x"346F" => data_out<= x"6E";
        when x"3470" => data_out<= x"29";
        when x"3471" => data_out<= x"0D";
        when x"3472" => data_out<= x"0A";
        when x"3473" => data_out<= x"00";
        when x"3474" => data_out<= x"43";
        when x"3475" => data_out<= x"41";
        when x"3476" => data_out<= x"54";
        when x"3477" => data_out<= x"20";
        when x"3478" => data_out<= x"66";
        when x"3479" => data_out<= x"69";
        when x"347A" => data_out<= x"6C";
        when x"347B" => data_out<= x"65";
        when x"347C" => data_out<= x"20";
        when x"347D" => data_out<= x"2D";
        when x"347E" => data_out<= x"20";
        when x"347F" => data_out<= x"56";
        when x"3480" => data_out<= x"65";
        when x"3481" => data_out<= x"72";
        when x"3482" => data_out<= x"20";
        when x"3483" => data_out<= x"63";
        when x"3484" => data_out<= x"6F";
        when x"3485" => data_out<= x"6E";
        when x"3486" => data_out<= x"74";
        when x"3487" => data_out<= x"65";
        when x"3488" => data_out<= x"6E";
        when x"3489" => data_out<= x"69";
        when x"348A" => data_out<= x"64";
        when x"348B" => data_out<= x"6F";
        when x"348C" => data_out<= x"20";
        when x"348D" => data_out<= x"68";
        when x"348E" => data_out<= x"65";
        when x"348F" => data_out<= x"78";
        when x"3490" => data_out<= x"0D";
        when x"3491" => data_out<= x"0A";
        when x"3492" => data_out<= x"00";
        when x"3493" => data_out<= x"44";
        when x"3494" => data_out<= x"65";
        when x"3495" => data_out<= x"62";
        when x"3496" => data_out<= x"65";
        when x"3497" => data_out<= x"20";
        when x"3498" => data_out<= x"74";
        when x"3499" => data_out<= x"65";
        when x"349A" => data_out<= x"72";
        when x"349B" => data_out<= x"6D";
        when x"349C" => data_out<= x"69";
        when x"349D" => data_out<= x"6E";
        when x"349E" => data_out<= x"61";
        when x"349F" => data_out<= x"72";
        when x"34A0" => data_out<= x"20";
        when x"34A1" => data_out<= x"63";
        when x"34A2" => data_out<= x"6F";
        when x"34A3" => data_out<= x"6E";
        when x"34A4" => data_out<= x"20";
        when x"34A5" => data_out<= x"52";
        when x"34A6" => data_out<= x"54";
        when x"34A7" => data_out<= x"53";
        when x"34A8" => data_out<= x"20";
        when x"34A9" => data_out<= x"28";
        when x"34AA" => data_out<= x"24";
        when x"34AB" => data_out<= x"36";
        when x"34AC" => data_out<= x"30";
        when x"34AD" => data_out<= x"29";
        when x"34AE" => data_out<= x"0D";
        when x"34AF" => data_out<= x"0A";
        when x"34B0" => data_out<= x"00";
        when x"34B1" => data_out<= x"53";
        when x"34B2" => data_out<= x"44";
        when x"34B3" => data_out<= x"20";
        when x"34B4" => data_out<= x"6E";
        when x"34B5" => data_out<= x"6F";
        when x"34B6" => data_out<= x"20";
        when x"34B7" => data_out<= x"6D";
        when x"34B8" => data_out<= x"6F";
        when x"34B9" => data_out<= x"6E";
        when x"34BA" => data_out<= x"74";
        when x"34BB" => data_out<= x"61";
        when x"34BC" => data_out<= x"64";
        when x"34BD" => data_out<= x"61";
        when x"34BE" => data_out<= x"2E";
        when x"34BF" => data_out<= x"20";
        when x"34C0" => data_out<= x"55";
        when x"34C1" => data_out<= x"73";
        when x"34C2" => data_out<= x"65";
        when x"34C3" => data_out<= x"20";
        when x"34C4" => data_out<= x"53";
        when x"34C5" => data_out<= x"44";
        when x"34C6" => data_out<= x"20";
        when x"34C7" => data_out<= x"70";
        when x"34C8" => data_out<= x"72";
        when x"34C9" => data_out<= x"69";
        when x"34CA" => data_out<= x"6D";
        when x"34CB" => data_out<= x"65";
        when x"34CC" => data_out<= x"72";
        when x"34CD" => data_out<= x"6F";
        when x"34CE" => data_out<= x"00";
        when x"34CF" => data_out<= x"44";
        when x"34D0" => data_out<= x"45";
        when x"34D1" => data_out<= x"4C";
        when x"34D2" => data_out<= x"20";
        when x"34D3" => data_out<= x"66";
        when x"34D4" => data_out<= x"69";
        when x"34D5" => data_out<= x"6C";
        when x"34D6" => data_out<= x"65";
        when x"34D7" => data_out<= x"20";
        when x"34D8" => data_out<= x"2D";
        when x"34D9" => data_out<= x"20";
        when x"34DA" => data_out<= x"45";
        when x"34DB" => data_out<= x"6C";
        when x"34DC" => data_out<= x"69";
        when x"34DD" => data_out<= x"6D";
        when x"34DE" => data_out<= x"69";
        when x"34DF" => data_out<= x"6E";
        when x"34E0" => data_out<= x"61";
        when x"34E1" => data_out<= x"72";
        when x"34E2" => data_out<= x"20";
        when x"34E3" => data_out<= x"61";
        when x"34E4" => data_out<= x"72";
        when x"34E5" => data_out<= x"63";
        when x"34E6" => data_out<= x"68";
        when x"34E7" => data_out<= x"69";
        when x"34E8" => data_out<= x"76";
        when x"34E9" => data_out<= x"6F";
        when x"34EA" => data_out<= x"0D";
        when x"34EB" => data_out<= x"0A";
        when x"34EC" => data_out<= x"00";
        when x"34ED" => data_out<= x"43";
        when x"34EE" => data_out<= x"6D";
        when x"34EF" => data_out<= x"64";
        when x"34F0" => data_out<= x"20";
        when x"34F1" => data_out<= x"64";
        when x"34F2" => data_out<= x"65";
        when x"34F3" => data_out<= x"73";
        when x"34F4" => data_out<= x"68";
        when x"34F5" => data_out<= x"61";
        when x"34F6" => data_out<= x"62";
        when x"34F7" => data_out<= x"69";
        when x"34F8" => data_out<= x"6C";
        when x"34F9" => data_out<= x"69";
        when x"34FA" => data_out<= x"74";
        when x"34FB" => data_out<= x"61";
        when x"34FC" => data_out<= x"64";
        when x"34FD" => data_out<= x"6F";
        when x"34FE" => data_out<= x"20";
        when x"34FF" => data_out<= x"70";
        when x"3500" => data_out<= x"2F";
        when x"3501" => data_out<= x"20";
        when x"3502" => data_out<= x"58";
        when x"3503" => data_out<= x"4D";
        when x"3504" => data_out<= x"4F";
        when x"3505" => data_out<= x"44";
        when x"3506" => data_out<= x"45";
        when x"3507" => data_out<= x"4D";
        when x"3508" => data_out<= x"0D";
        when x"3509" => data_out<= x"0A";
        when x"350A" => data_out<= x"00";
        when x"350B" => data_out<= x"45";
        when x"350C" => data_out<= x"6A";
        when x"350D" => data_out<= x"3A";
        when x"350E" => data_out<= x"20";
        when x"350F" => data_out<= x"53";
        when x"3510" => data_out<= x"41";
        when x"3511" => data_out<= x"56";
        when x"3512" => data_out<= x"45";
        when x"3513" => data_out<= x"20";
        when x"3514" => data_out<= x"50";
        when x"3515" => data_out<= x"52";
        when x"3516" => data_out<= x"4F";
        when x"3517" => data_out<= x"47";
        when x"3518" => data_out<= x"2E";
        when x"3519" => data_out<= x"42";
        when x"351A" => data_out<= x"49";
        when x"351B" => data_out<= x"4E";
        when x"351C" => data_out<= x"20";
        when x"351D" => data_out<= x"30";
        when x"351E" => data_out<= x"32";
        when x"351F" => data_out<= x"30";
        when x"3520" => data_out<= x"30";
        when x"3521" => data_out<= x"20";
        when x"3522" => data_out<= x"31";
        when x"3523" => data_out<= x"30";
        when x"3524" => data_out<= x"30";
        when x"3525" => data_out<= x"0D";
        when x"3526" => data_out<= x"0A";
        when x"3527" => data_out<= x"00";
        when x"3528" => data_out<= x"57";
        when x"3529" => data_out<= x"20";
        when x"352A" => data_out<= x"61";
        when x"352B" => data_out<= x"64";
        when x"352C" => data_out<= x"64";
        when x"352D" => data_out<= x"72";
        when x"352E" => data_out<= x"20";
        when x"352F" => data_out<= x"76";
        when x"3530" => data_out<= x"61";
        when x"3531" => data_out<= x"6C";
        when x"3532" => data_out<= x"20";
        when x"3533" => data_out<= x"2D";
        when x"3534" => data_out<= x"20";
        when x"3535" => data_out<= x"45";
        when x"3536" => data_out<= x"73";
        when x"3537" => data_out<= x"63";
        when x"3538" => data_out<= x"72";
        when x"3539" => data_out<= x"69";
        when x"353A" => data_out<= x"62";
        when x"353B" => data_out<= x"69";
        when x"353C" => data_out<= x"72";
        when x"353D" => data_out<= x"20";
        when x"353E" => data_out<= x"62";
        when x"353F" => data_out<= x"79";
        when x"3540" => data_out<= x"74";
        when x"3541" => data_out<= x"65";
        when x"3542" => data_out<= x"0D";
        when x"3543" => data_out<= x"0A";
        when x"3544" => data_out<= x"00";
        when x"3545" => data_out<= x"52";
        when x"3546" => data_out<= x"20";
        when x"3547" => data_out<= x"5B";
        when x"3548" => data_out<= x"61";
        when x"3549" => data_out<= x"64";
        when x"354A" => data_out<= x"64";
        when x"354B" => data_out<= x"72";
        when x"354C" => data_out<= x"5D";
        when x"354D" => data_out<= x"20";
        when x"354E" => data_out<= x"20";
        when x"354F" => data_out<= x"20";
        when x"3550" => data_out<= x"52";
        when x"3551" => data_out<= x"75";
        when x"3552" => data_out<= x"6E";
        when x"3553" => data_out<= x"20";
        when x"3554" => data_out<= x"28";
        when x"3555" => data_out<= x"64";
        when x"3556" => data_out<= x"65";
        when x"3557" => data_out<= x"66";
        when x"3558" => data_out<= x"20";
        when x"3559" => data_out<= x"24";
        when x"355A" => data_out<= x"30";
        when x"355B" => data_out<= x"38";
        when x"355C" => data_out<= x"30";
        when x"355D" => data_out<= x"30";
        when x"355E" => data_out<= x"29";
        when x"355F" => data_out<= x"0D";
        when x"3560" => data_out<= x"0A";
        when x"3561" => data_out<= x"00";
        when x"3562" => data_out<= x"43";
        when x"3563" => data_out<= x"6F";
        when x"3564" => data_out<= x"6D";
        when x"3565" => data_out<= x"61";
        when x"3566" => data_out<= x"6E";
        when x"3567" => data_out<= x"64";
        when x"3568" => data_out<= x"6F";
        when x"3569" => data_out<= x"20";
        when x"356A" => data_out<= x"64";
        when x"356B" => data_out<= x"65";
        when x"356C" => data_out<= x"73";
        when x"356D" => data_out<= x"63";
        when x"356E" => data_out<= x"6F";
        when x"356F" => data_out<= x"6E";
        when x"3570" => data_out<= x"6F";
        when x"3571" => data_out<= x"63";
        when x"3572" => data_out<= x"69";
        when x"3573" => data_out<= x"64";
        when x"3574" => data_out<= x"6F";
        when x"3575" => data_out<= x"2E";
        when x"3576" => data_out<= x"20";
        when x"3577" => data_out<= x"48";
        when x"3578" => data_out<= x"3D";
        when x"3579" => data_out<= x"61";
        when x"357A" => data_out<= x"79";
        when x"357B" => data_out<= x"75";
        when x"357C" => data_out<= x"64";
        when x"357D" => data_out<= x"61";
        when x"357E" => data_out<= x"00";
        when x"357F" => data_out<= x"20";
        when x"3580" => data_out<= x"20";
        when x"3581" => data_out<= x"53";
        when x"3582" => data_out<= x"69";
        when x"3583" => data_out<= x"6E";
        when x"3584" => data_out<= x"20";
        when x"3585" => data_out<= x"46";
        when x"3586" => data_out<= x"53";
        when x"3587" => data_out<= x"2E";
        when x"3588" => data_out<= x"20";
        when x"3589" => data_out<= x"46";
        when x"358A" => data_out<= x"6F";
        when x"358B" => data_out<= x"72";
        when x"358C" => data_out<= x"6D";
        when x"358D" => data_out<= x"61";
        when x"358E" => data_out<= x"74";
        when x"358F" => data_out<= x"65";
        when x"3590" => data_out<= x"61";
        when x"3591" => data_out<= x"72";
        when x"3592" => data_out<= x"3F";
        when x"3593" => data_out<= x"20";
        when x"3594" => data_out<= x"28";
        when x"3595" => data_out<= x"53";
        when x"3596" => data_out<= x"2F";
        when x"3597" => data_out<= x"4E";
        when x"3598" => data_out<= x"29";
        when x"3599" => data_out<= x"3A";
        when x"359A" => data_out<= x"20";
        when x"359B" => data_out<= x"00";
        when x"359C" => data_out<= x"45";
        when x"359D" => data_out<= x"73";
        when x"359E" => data_out<= x"63";
        when x"359F" => data_out<= x"72";
        when x"35A0" => data_out<= x"69";
        when x"35A1" => data_out<= x"62";
        when x"35A2" => data_out<= x"65";
        when x"35A3" => data_out<= x"20";
        when x"35A4" => data_out<= x"62";
        when x"35A5" => data_out<= x"79";
        when x"35A6" => data_out<= x"74";
        when x"35A7" => data_out<= x"65";
        when x"35A8" => data_out<= x"73";
        when x"35A9" => data_out<= x"2C";
        when x"35AA" => data_out<= x"20";
        when x"35AB" => data_out<= x"27";
        when x"35AC" => data_out<= x"2E";
        when x"35AD" => data_out<= x"27";
        when x"35AE" => data_out<= x"20";
        when x"35AF" => data_out<= x"74";
        when x"35B0" => data_out<= x"65";
        when x"35B1" => data_out<= x"72";
        when x"35B2" => data_out<= x"6D";
        when x"35B3" => data_out<= x"69";
        when x"35B4" => data_out<= x"6E";
        when x"35B5" => data_out<= x"61";
        when x"35B6" => data_out<= x"0D";
        when x"35B7" => data_out<= x"0A";
        when x"35B8" => data_out<= x"00";
        when x"35B9" => data_out<= x"4D";
        when x"35BA" => data_out<= x"20";
        when x"35BB" => data_out<= x"61";
        when x"35BC" => data_out<= x"64";
        when x"35BD" => data_out<= x"64";
        when x"35BE" => data_out<= x"72";
        when x"35BF" => data_out<= x"20";
        when x"35C0" => data_out<= x"5B";
        when x"35C1" => data_out<= x"6E";
        when x"35C2" => data_out<= x"5D";
        when x"35C3" => data_out<= x"20";
        when x"35C4" => data_out<= x"2D";
        when x"35C5" => data_out<= x"20";
        when x"35C6" => data_out<= x"44";
        when x"35C7" => data_out<= x"65";
        when x"35C8" => data_out<= x"73";
        when x"35C9" => data_out<= x"65";
        when x"35CA" => data_out<= x"6E";
        when x"35CB" => data_out<= x"73";
        when x"35CC" => data_out<= x"61";
        when x"35CD" => data_out<= x"6D";
        when x"35CE" => data_out<= x"62";
        when x"35CF" => data_out<= x"6C";
        when x"35D0" => data_out<= x"61";
        when x"35D1" => data_out<= x"72";
        when x"35D2" => data_out<= x"0D";
        when x"35D3" => data_out<= x"0A";
        when x"35D4" => data_out<= x"00";
        when x"35D5" => data_out<= x"42";
        when x"35D6" => data_out<= x"4F";
        when x"35D7" => data_out<= x"52";
        when x"35D8" => data_out<= x"52";
        when x"35D9" => data_out<= x"41";
        when x"35DA" => data_out<= x"20";
        when x"35DB" => data_out<= x"74";
        when x"35DC" => data_out<= x"6F";
        when x"35DD" => data_out<= x"64";
        when x"35DE" => data_out<= x"6F";
        when x"35DF" => data_out<= x"73";
        when x"35E0" => data_out<= x"20";
        when x"35E1" => data_out<= x"6C";
        when x"35E2" => data_out<= x"6F";
        when x"35E3" => data_out<= x"73";
        when x"35E4" => data_out<= x"20";
        when x"35E5" => data_out<= x"61";
        when x"35E6" => data_out<= x"72";
        when x"35E7" => data_out<= x"63";
        when x"35E8" => data_out<= x"68";
        when x"35E9" => data_out<= x"69";
        when x"35EA" => data_out<= x"76";
        when x"35EB" => data_out<= x"6F";
        when x"35EC" => data_out<= x"73";
        when x"35ED" => data_out<= x"21";
        when x"35EE" => data_out<= x"0D";
        when x"35EF" => data_out<= x"0A";
        when x"35F0" => data_out<= x"00";
        when x"35F1" => data_out<= x"6E";
        when x"35F2" => data_out<= x"3D";
        when x"35F3" => data_out<= x"69";
        when x"35F4" => data_out<= x"6E";
        when x"35F5" => data_out<= x"73";
        when x"35F6" => data_out<= x"74";
        when x"35F7" => data_out<= x"72";
        when x"35F8" => data_out<= x"75";
        when x"35F9" => data_out<= x"63";
        when x"35FA" => data_out<= x"63";
        when x"35FB" => data_out<= x"69";
        when x"35FC" => data_out<= x"6F";
        when x"35FD" => data_out<= x"6E";
        when x"35FE" => data_out<= x"65";
        when x"35FF" => data_out<= x"73";
        when x"3600" => data_out<= x"20";
        when x"3601" => data_out<= x"28";
        when x"3602" => data_out<= x"64";
        when x"3603" => data_out<= x"65";
        when x"3604" => data_out<= x"66";
        when x"3605" => data_out<= x"20";
        when x"3606" => data_out<= x"31";
        when x"3607" => data_out<= x"36";
        when x"3608" => data_out<= x"29";
        when x"3609" => data_out<= x"0D";
        when x"360A" => data_out<= x"0A";
        when x"360B" => data_out<= x"00";
        when x"360C" => data_out<= x"53";
        when x"360D" => data_out<= x"44";
        when x"360E" => data_out<= x"20";
        when x"360F" => data_out<= x"2D";
        when x"3610" => data_out<= x"20";
        when x"3611" => data_out<= x"49";
        when x"3612" => data_out<= x"6E";
        when x"3613" => data_out<= x"69";
        when x"3614" => data_out<= x"63";
        when x"3615" => data_out<= x"69";
        when x"3616" => data_out<= x"61";
        when x"3617" => data_out<= x"6C";
        when x"3618" => data_out<= x"69";
        when x"3619" => data_out<= x"7A";
        when x"361A" => data_out<= x"61";
        when x"361B" => data_out<= x"72";
        when x"361C" => data_out<= x"20";
        when x"361D" => data_out<= x"53";
        when x"361E" => data_out<= x"44";
        when x"361F" => data_out<= x"20";
        when x"3620" => data_out<= x"43";
        when x"3621" => data_out<= x"61";
        when x"3622" => data_out<= x"72";
        when x"3623" => data_out<= x"64";
        when x"3624" => data_out<= x"0D";
        when x"3625" => data_out<= x"0A";
        when x"3626" => data_out<= x"00";
        when x"3627" => data_out<= x"20";
        when x"3628" => data_out<= x"20";
        when x"3629" => data_out<= x"4D";
        when x"362A" => data_out<= x"4F";
        when x"362B" => data_out<= x"4E";
        when x"362C" => data_out<= x"49";
        when x"362D" => data_out<= x"54";
        when x"362E" => data_out<= x"4F";
        when x"362F" => data_out<= x"52";
        when x"3630" => data_out<= x"20";
        when x"3631" => data_out<= x"36";
        when x"3632" => data_out<= x"35";
        when x"3633" => data_out<= x"30";
        when x"3634" => data_out<= x"32";
        when x"3635" => data_out<= x"20";
        when x"3636" => data_out<= x"76";
        when x"3637" => data_out<= x"32";
        when x"3638" => data_out<= x"2E";
        when x"3639" => data_out<= x"33";
        when x"363A" => data_out<= x"2E";
        when x"363B" => data_out<= x"30";
        when x"363C" => data_out<= x"20";
        when x"363D" => data_out<= x"2B";
        when x"363E" => data_out<= x"20";
        when x"363F" => data_out<= x"53";
        when x"3640" => data_out<= x"44";
        when x"3641" => data_out<= x"00";
        when x"3642" => data_out<= x"20";
        when x"3643" => data_out<= x"20";
        when x"3644" => data_out<= x"54";
        when x"3645" => data_out<= x"61";
        when x"3646" => data_out<= x"6E";
        when x"3647" => data_out<= x"67";
        when x"3648" => data_out<= x"20";
        when x"3649" => data_out<= x"4E";
        when x"364A" => data_out<= x"61";
        when x"364B" => data_out<= x"6E";
        when x"364C" => data_out<= x"6F";
        when x"364D" => data_out<= x"20";
        when x"364E" => data_out<= x"39";
        when x"364F" => data_out<= x"4B";
        when x"3650" => data_out<= x"20";
        when x"3651" => data_out<= x"40";
        when x"3652" => data_out<= x"20";
        when x"3653" => data_out<= x"33";
        when x"3654" => data_out<= x"2E";
        when x"3655" => data_out<= x"33";
        when x"3656" => data_out<= x"37";
        when x"3657" => data_out<= x"35";
        when x"3658" => data_out<= x"20";
        when x"3659" => data_out<= x"4D";
        when x"365A" => data_out<= x"48";
        when x"365B" => data_out<= x"7A";
        when x"365C" => data_out<= x"00";
        when x"365D" => data_out<= x"45";
        when x"365E" => data_out<= x"6A";
        when x"365F" => data_out<= x"3A";
        when x"3660" => data_out<= x"20";
        when x"3661" => data_out<= x"57";
        when x"3662" => data_out<= x"20";
        when x"3663" => data_out<= x"30";
        when x"3664" => data_out<= x"32";
        when x"3665" => data_out<= x"30";
        when x"3666" => data_out<= x"30";
        when x"3667" => data_out<= x"20";
        when x"3668" => data_out<= x"46";
        when x"3669" => data_out<= x"46";
        when x"366A" => data_out<= x"2C";
        when x"366B" => data_out<= x"20";
        when x"366C" => data_out<= x"57";
        when x"366D" => data_out<= x"20";
        when x"366E" => data_out<= x"43";
        when x"366F" => data_out<= x"30";
        when x"3670" => data_out<= x"30";
        when x"3671" => data_out<= x"31";
        when x"3672" => data_out<= x"20";
        when x"3673" => data_out<= x"33";
        when x"3674" => data_out<= x"46";
        when x"3675" => data_out<= x"0D";
        when x"3676" => data_out<= x"0A";
        when x"3677" => data_out<= x"00";
        when x"3678" => data_out<= x"49";
        when x"3679" => data_out<= x"20";
        when x"367A" => data_out<= x"20";
        when x"367B" => data_out<= x"20";
        when x"367C" => data_out<= x"20";
        when x"367D" => data_out<= x"20";
        when x"367E" => data_out<= x"20";
        when x"367F" => data_out<= x"20";
        when x"3680" => data_out<= x"20";
        when x"3681" => data_out<= x"20";
        when x"3682" => data_out<= x"20";
        when x"3683" => data_out<= x"49";
        when x"3684" => data_out<= x"6E";
        when x"3685" => data_out<= x"66";
        when x"3686" => data_out<= x"6F";
        when x"3687" => data_out<= x"20";
        when x"3688" => data_out<= x"6D";
        when x"3689" => data_out<= x"65";
        when x"368A" => data_out<= x"6D";
        when x"368B" => data_out<= x"6F";
        when x"368C" => data_out<= x"72";
        when x"368D" => data_out<= x"69";
        when x"368E" => data_out<= x"61";
        when x"368F" => data_out<= x"0D";
        when x"3690" => data_out<= x"0A";
        when x"3691" => data_out<= x"00";
        when x"3692" => data_out<= x"55";
        when x"3693" => data_out<= x"73";
        when x"3694" => data_out<= x"6F";
        when x"3695" => data_out<= x"3A";
        when x"3696" => data_out<= x"20";
        when x"3697" => data_out<= x"53";
        when x"3698" => data_out<= x"41";
        when x"3699" => data_out<= x"56";
        when x"369A" => data_out<= x"45";
        when x"369B" => data_out<= x"20";
        when x"369C" => data_out<= x"6E";
        when x"369D" => data_out<= x"6F";
        when x"369E" => data_out<= x"6D";
        when x"369F" => data_out<= x"62";
        when x"36A0" => data_out<= x"72";
        when x"36A1" => data_out<= x"65";
        when x"36A2" => data_out<= x"20";
        when x"36A3" => data_out<= x"61";
        when x"36A4" => data_out<= x"64";
        when x"36A5" => data_out<= x"64";
        when x"36A6" => data_out<= x"72";
        when x"36A7" => data_out<= x"20";
        when x"36A8" => data_out<= x"6C";
        when x"36A9" => data_out<= x"65";
        when x"36AA" => data_out<= x"6E";
        when x"36AB" => data_out<= x"00";
        when x"36AC" => data_out<= x"53";
        when x"36AD" => data_out<= x"44";
        when x"36AE" => data_out<= x"46";
        when x"36AF" => data_out<= x"4F";
        when x"36B0" => data_out<= x"52";
        when x"36B1" => data_out<= x"4D";
        when x"36B2" => data_out<= x"41";
        when x"36B3" => data_out<= x"54";
        when x"36B4" => data_out<= x"20";
        when x"36B5" => data_out<= x"2D";
        when x"36B6" => data_out<= x"20";
        when x"36B7" => data_out<= x"46";
        when x"36B8" => data_out<= x"6F";
        when x"36B9" => data_out<= x"72";
        when x"36BA" => data_out<= x"6D";
        when x"36BB" => data_out<= x"61";
        when x"36BC" => data_out<= x"74";
        when x"36BD" => data_out<= x"65";
        when x"36BE" => data_out<= x"61";
        when x"36BF" => data_out<= x"72";
        when x"36C0" => data_out<= x"20";
        when x"36C1" => data_out<= x"53";
        when x"36C2" => data_out<= x"44";
        when x"36C3" => data_out<= x"0D";
        when x"36C4" => data_out<= x"0A";
        when x"36C5" => data_out<= x"00";
        when x"36C6" => data_out<= x"4D";
        when x"36C7" => data_out<= x"75";
        when x"36C8" => data_out<= x"65";
        when x"36C9" => data_out<= x"73";
        when x"36CA" => data_out<= x"74";
        when x"36CB" => data_out<= x"72";
        when x"36CC" => data_out<= x"61";
        when x"36CD" => data_out<= x"20";
        when x"36CE" => data_out<= x"6E";
        when x"36CF" => data_out<= x"6F";
        when x"36D0" => data_out<= x"6D";
        when x"36D1" => data_out<= x"62";
        when x"36D2" => data_out<= x"72";
        when x"36D3" => data_out<= x"65";
        when x"36D4" => data_out<= x"20";
        when x"36D5" => data_out<= x"79";
        when x"36D6" => data_out<= x"20";
        when x"36D7" => data_out<= x"74";
        when x"36D8" => data_out<= x"61";
        when x"36D9" => data_out<= x"6D";
        when x"36DA" => data_out<= x"61";
        when x"36DB" => data_out<= x"6E";
        when x"36DC" => data_out<= x"6F";
        when x"36DD" => data_out<= x"0D";
        when x"36DE" => data_out<= x"0A";
        when x"36DF" => data_out<= x"00";
        when x"36E0" => data_out<= x"52";
        when x"36E1" => data_out<= x"41";
        when x"36E2" => data_out<= x"4D";
        when x"36E3" => data_out<= x"3A";
        when x"36E4" => data_out<= x"20";
        when x"36E5" => data_out<= x"20";
        when x"36E6" => data_out<= x"20";
        when x"36E7" => data_out<= x"20";
        when x"36E8" => data_out<= x"20";
        when x"36E9" => data_out<= x"20";
        when x"36EA" => data_out<= x"20";
        when x"36EB" => data_out<= x"20";
        when x"36EC" => data_out<= x"24";
        when x"36ED" => data_out<= x"30";
        when x"36EE" => data_out<= x"31";
        when x"36EF" => data_out<= x"30";
        when x"36F0" => data_out<= x"30";
        when x"36F1" => data_out<= x"2D";
        when x"36F2" => data_out<= x"24";
        when x"36F3" => data_out<= x"33";
        when x"36F4" => data_out<= x"44";
        when x"36F5" => data_out<= x"46";
        when x"36F6" => data_out<= x"46";
        when x"36F7" => data_out<= x"20";
        when x"36F8" => data_out<= x"28";
        when x"36F9" => data_out<= x"00";
        when x"36FA" => data_out<= x"5A";
        when x"36FB" => data_out<= x"65";
        when x"36FC" => data_out<= x"72";
        when x"36FD" => data_out<= x"6F";
        when x"36FE" => data_out<= x"20";
        when x"36FF" => data_out<= x"50";
        when x"3700" => data_out<= x"61";
        when x"3701" => data_out<= x"67";
        when x"3702" => data_out<= x"65";
        when x"3703" => data_out<= x"3A";
        when x"3704" => data_out<= x"20";
        when x"3705" => data_out<= x"20";
        when x"3706" => data_out<= x"24";
        when x"3707" => data_out<= x"30";
        when x"3708" => data_out<= x"30";
        when x"3709" => data_out<= x"30";
        when x"370A" => data_out<= x"32";
        when x"370B" => data_out<= x"2D";
        when x"370C" => data_out<= x"24";
        when x"370D" => data_out<= x"30";
        when x"370E" => data_out<= x"30";
        when x"370F" => data_out<= x"46";
        when x"3710" => data_out<= x"46";
        when x"3711" => data_out<= x"20";
        when x"3712" => data_out<= x"28";
        when x"3713" => data_out<= x"00";
        when x"3714" => data_out<= x"43";
        when x"3715" => data_out<= x"61";
        when x"3716" => data_out<= x"72";
        when x"3717" => data_out<= x"67";
        when x"3718" => data_out<= x"61";
        when x"3719" => data_out<= x"20";
        when x"371A" => data_out<= x"61";
        when x"371B" => data_out<= x"72";
        when x"371C" => data_out<= x"63";
        when x"371D" => data_out<= x"68";
        when x"371E" => data_out<= x"69";
        when x"371F" => data_out<= x"76";
        when x"3720" => data_out<= x"6F";
        when x"3721" => data_out<= x"20";
        when x"3722" => data_out<= x"61";
        when x"3723" => data_out<= x"20";
        when x"3724" => data_out<= x"6D";
        when x"3725" => data_out<= x"65";
        when x"3726" => data_out<= x"6D";
        when x"3727" => data_out<= x"6F";
        when x"3728" => data_out<= x"72";
        when x"3729" => data_out<= x"69";
        when x"372A" => data_out<= x"61";
        when x"372B" => data_out<= x"0D";
        when x"372C" => data_out<= x"0A";
        when x"372D" => data_out<= x"00";
        when x"372E" => data_out<= x"53";
        when x"372F" => data_out<= x"74";
        when x"3730" => data_out<= x"61";
        when x"3731" => data_out<= x"63";
        when x"3732" => data_out<= x"6B";
        when x"3733" => data_out<= x"3A";
        when x"3734" => data_out<= x"20";
        when x"3735" => data_out<= x"20";
        when x"3736" => data_out<= x"20";
        when x"3737" => data_out<= x"20";
        when x"3738" => data_out<= x"20";
        when x"3739" => data_out<= x"20";
        when x"373A" => data_out<= x"24";
        when x"373B" => data_out<= x"33";
        when x"373C" => data_out<= x"45";
        when x"373D" => data_out<= x"30";
        when x"373E" => data_out<= x"30";
        when x"373F" => data_out<= x"2D";
        when x"3740" => data_out<= x"24";
        when x"3741" => data_out<= x"33";
        when x"3742" => data_out<= x"46";
        when x"3743" => data_out<= x"46";
        when x"3744" => data_out<= x"46";
        when x"3745" => data_out<= x"20";
        when x"3746" => data_out<= x"28";
        when x"3747" => data_out<= x"00";
        when x"3748" => data_out<= x"4C";
        when x"3749" => data_out<= x"53";
        when x"374A" => data_out<= x"20";
        when x"374B" => data_out<= x"2D";
        when x"374C" => data_out<= x"20";
        when x"374D" => data_out<= x"4C";
        when x"374E" => data_out<= x"69";
        when x"374F" => data_out<= x"73";
        when x"3750" => data_out<= x"74";
        when x"3751" => data_out<= x"61";
        when x"3752" => data_out<= x"72";
        when x"3753" => data_out<= x"20";
        when x"3754" => data_out<= x"61";
        when x"3755" => data_out<= x"72";
        when x"3756" => data_out<= x"63";
        when x"3757" => data_out<= x"68";
        when x"3758" => data_out<= x"69";
        when x"3759" => data_out<= x"76";
        when x"375A" => data_out<= x"6F";
        when x"375B" => data_out<= x"73";
        when x"375C" => data_out<= x"20";
        when x"375D" => data_out<= x"53";
        when x"375E" => data_out<= x"44";
        when x"375F" => data_out<= x"0D";
        when x"3760" => data_out<= x"0A";
        when x"3761" => data_out<= x"00";
        when x"3762" => data_out<= x"4D";
        when x"3763" => data_out<= x"20";
        when x"3764" => data_out<= x"61";
        when x"3765" => data_out<= x"64";
        when x"3766" => data_out<= x"64";
        when x"3767" => data_out<= x"72";
        when x"3768" => data_out<= x"20";
        when x"3769" => data_out<= x"5B";
        when x"376A" => data_out<= x"6E";
        when x"376B" => data_out<= x"5D";
        when x"376C" => data_out<= x"20";
        when x"376D" => data_out<= x"44";
        when x"376E" => data_out<= x"65";
        when x"376F" => data_out<= x"73";
        when x"3770" => data_out<= x"65";
        when x"3771" => data_out<= x"6E";
        when x"3772" => data_out<= x"73";
        when x"3773" => data_out<= x"61";
        when x"3774" => data_out<= x"6D";
        when x"3775" => data_out<= x"62";
        when x"3776" => data_out<= x"6C";
        when x"3777" => data_out<= x"61";
        when x"3778" => data_out<= x"72";
        when x"3779" => data_out<= x"0D";
        when x"377A" => data_out<= x"0A";
        when x"377B" => data_out<= x"00";
        when x"377C" => data_out<= x"49";
        when x"377D" => data_out<= x"6E";
        when x"377E" => data_out<= x"69";
        when x"377F" => data_out<= x"63";
        when x"3780" => data_out<= x"69";
        when x"3781" => data_out<= x"61";
        when x"3782" => data_out<= x"6C";
        when x"3783" => data_out<= x"69";
        when x"3784" => data_out<= x"7A";
        when x"3785" => data_out<= x"61";
        when x"3786" => data_out<= x"6E";
        when x"3787" => data_out<= x"64";
        when x"3788" => data_out<= x"6F";
        when x"3789" => data_out<= x"20";
        when x"378A" => data_out<= x"53";
        when x"378B" => data_out<= x"44";
        when x"378C" => data_out<= x"20";
        when x"378D" => data_out<= x"43";
        when x"378E" => data_out<= x"61";
        when x"378F" => data_out<= x"72";
        when x"3790" => data_out<= x"64";
        when x"3791" => data_out<= x"2E";
        when x"3792" => data_out<= x"2E";
        when x"3793" => data_out<= x"2E";
        when x"3794" => data_out<= x"00";
        when x"3795" => data_out<= x"4D";
        when x"3796" => data_out<= x"6F";
        when x"3797" => data_out<= x"6E";
        when x"3798" => data_out<= x"69";
        when x"3799" => data_out<= x"74";
        when x"379A" => data_out<= x"6F";
        when x"379B" => data_out<= x"72";
        when x"379C" => data_out<= x"20";
        when x"379D" => data_out<= x"42";
        when x"379E" => data_out<= x"53";
        when x"379F" => data_out<= x"53";
        when x"37A0" => data_out<= x"3A";
        when x"37A1" => data_out<= x"20";
        when x"37A2" => data_out<= x"24";
        when x"37A3" => data_out<= x"30";
        when x"37A4" => data_out<= x"32";
        when x"37A5" => data_out<= x"30";
        when x"37A6" => data_out<= x"30";
        when x"37A7" => data_out<= x"2D";
        when x"37A8" => data_out<= x"24";
        when x"37A9" => data_out<= x"30";
        when x"37AA" => data_out<= x"37";
        when x"37AB" => data_out<= x"46";
        when x"37AC" => data_out<= x"46";
        when x"37AD" => data_out<= x"00";
        when x"37AE" => data_out<= x"55";
        when x"37AF" => data_out<= x"73";
        when x"37B0" => data_out<= x"6F";
        when x"37B1" => data_out<= x"3A";
        when x"37B2" => data_out<= x"20";
        when x"37B3" => data_out<= x"4C";
        when x"37B4" => data_out<= x"4F";
        when x"37B5" => data_out<= x"41";
        when x"37B6" => data_out<= x"44";
        when x"37B7" => data_out<= x"20";
        when x"37B8" => data_out<= x"6E";
        when x"37B9" => data_out<= x"6F";
        when x"37BA" => data_out<= x"6D";
        when x"37BB" => data_out<= x"62";
        when x"37BC" => data_out<= x"72";
        when x"37BD" => data_out<= x"65";
        when x"37BE" => data_out<= x"20";
        when x"37BF" => data_out<= x"5B";
        when x"37C0" => data_out<= x"61";
        when x"37C1" => data_out<= x"64";
        when x"37C2" => data_out<= x"64";
        when x"37C3" => data_out<= x"72";
        when x"37C4" => data_out<= x"5D";
        when x"37C5" => data_out<= x"00";
        when x"37C6" => data_out<= x"49";
        when x"37C7" => data_out<= x"2F";
        when x"37C8" => data_out<= x"4F";
        when x"37C9" => data_out<= x"3A";
        when x"37CA" => data_out<= x"20";
        when x"37CB" => data_out<= x"20";
        when x"37CC" => data_out<= x"20";
        when x"37CD" => data_out<= x"20";
        when x"37CE" => data_out<= x"20";
        when x"37CF" => data_out<= x"20";
        when x"37D0" => data_out<= x"20";
        when x"37D1" => data_out<= x"20";
        when x"37D2" => data_out<= x"24";
        when x"37D3" => data_out<= x"43";
        when x"37D4" => data_out<= x"30";
        when x"37D5" => data_out<= x"30";
        when x"37D6" => data_out<= x"30";
        when x"37D7" => data_out<= x"2D";
        when x"37D8" => data_out<= x"24";
        when x"37D9" => data_out<= x"43";
        when x"37DA" => data_out<= x"30";
        when x"37DB" => data_out<= x"46";
        when x"37DC" => data_out<= x"46";
        when x"37DD" => data_out<= x"00";
        when x"37DE" => data_out<= x"45";
        when x"37DF" => data_out<= x"6A";
        when x"37E0" => data_out<= x"3A";
        when x"37E1" => data_out<= x"20";
        when x"37E2" => data_out<= x"4D";
        when x"37E3" => data_out<= x"20";
        when x"37E4" => data_out<= x"30";
        when x"37E5" => data_out<= x"32";
        when x"37E6" => data_out<= x"30";
        when x"37E7" => data_out<= x"30";
        when x"37E8" => data_out<= x"2C";
        when x"37E9" => data_out<= x"20";
        when x"37EA" => data_out<= x"4D";
        when x"37EB" => data_out<= x"20";
        when x"37EC" => data_out<= x"38";
        when x"37ED" => data_out<= x"30";
        when x"37EE" => data_out<= x"30";
        when x"37EF" => data_out<= x"30";
        when x"37F0" => data_out<= x"20";
        when x"37F1" => data_out<= x"32";
        when x"37F2" => data_out<= x"30";
        when x"37F3" => data_out<= x"0D";
        when x"37F4" => data_out<= x"0A";
        when x"37F5" => data_out<= x"00";
        when x"37F6" => data_out<= x"49";
        when x"37F7" => data_out<= x"20";
        when x"37F8" => data_out<= x"2D";
        when x"37F9" => data_out<= x"20";
        when x"37FA" => data_out<= x"49";
        when x"37FB" => data_out<= x"6E";
        when x"37FC" => data_out<= x"66";
        when x"37FD" => data_out<= x"6F";
        when x"37FE" => data_out<= x"20";
        when x"37FF" => data_out<= x"6D";
        when x"3800" => data_out<= x"61";
        when x"3801" => data_out<= x"70";
        when x"3802" => data_out<= x"61";
        when x"3803" => data_out<= x"20";
        when x"3804" => data_out<= x"6D";
        when x"3805" => data_out<= x"65";
        when x"3806" => data_out<= x"6D";
        when x"3807" => data_out<= x"6F";
        when x"3808" => data_out<= x"72";
        when x"3809" => data_out<= x"69";
        when x"380A" => data_out<= x"61";
        when x"380B" => data_out<= x"0D";
        when x"380C" => data_out<= x"0A";
        when x"380D" => data_out<= x"00";
        when x"380E" => data_out<= x"51";
        when x"380F" => data_out<= x"20";
        when x"3810" => data_out<= x"2D";
        when x"3811" => data_out<= x"20";
        when x"3812" => data_out<= x"53";
        when x"3813" => data_out<= x"61";
        when x"3814" => data_out<= x"6C";
        when x"3815" => data_out<= x"69";
        when x"3816" => data_out<= x"72";
        when x"3817" => data_out<= x"20";
        when x"3818" => data_out<= x"64";
        when x"3819" => data_out<= x"65";
        when x"381A" => data_out<= x"6C";
        when x"381B" => data_out<= x"20";
        when x"381C" => data_out<= x"6D";
        when x"381D" => data_out<= x"6F";
        when x"381E" => data_out<= x"6E";
        when x"381F" => data_out<= x"69";
        when x"3820" => data_out<= x"74";
        when x"3821" => data_out<= x"6F";
        when x"3822" => data_out<= x"72";
        when x"3823" => data_out<= x"0D";
        when x"3824" => data_out<= x"0A";
        when x"3825" => data_out<= x"00";
        when x"3826" => data_out<= x"45";
        when x"3827" => data_out<= x"6A";
        when x"3828" => data_out<= x"3A";
        when x"3829" => data_out<= x"20";
        when x"382A" => data_out<= x"52";
        when x"382B" => data_out<= x"2C";
        when x"382C" => data_out<= x"20";
        when x"382D" => data_out<= x"52";
        when x"382E" => data_out<= x"20";
        when x"382F" => data_out<= x"30";
        when x"3830" => data_out<= x"38";
        when x"3831" => data_out<= x"30";
        when x"3832" => data_out<= x"30";
        when x"3833" => data_out<= x"2C";
        when x"3834" => data_out<= x"20";
        when x"3835" => data_out<= x"52";
        when x"3836" => data_out<= x"20";
        when x"3837" => data_out<= x"31";
        when x"3838" => data_out<= x"30";
        when x"3839" => data_out<= x"30";
        when x"383A" => data_out<= x"30";
        when x"383B" => data_out<= x"0D";
        when x"383C" => data_out<= x"0A";
        when x"383D" => data_out<= x"00";
        when x"383E" => data_out<= x"53";
        when x"383F" => data_out<= x"61";
        when x"3840" => data_out<= x"6C";
        when x"3841" => data_out<= x"69";
        when x"3842" => data_out<= x"65";
        when x"3843" => data_out<= x"6E";
        when x"3844" => data_out<= x"64";
        when x"3845" => data_out<= x"6F";
        when x"3846" => data_out<= x"20";
        when x"3847" => data_out<= x"64";
        when x"3848" => data_out<= x"65";
        when x"3849" => data_out<= x"6C";
        when x"384A" => data_out<= x"20";
        when x"384B" => data_out<= x"6D";
        when x"384C" => data_out<= x"6F";
        when x"384D" => data_out<= x"6E";
        when x"384E" => data_out<= x"69";
        when x"384F" => data_out<= x"74";
        when x"3850" => data_out<= x"6F";
        when x"3851" => data_out<= x"72";
        when x"3852" => data_out<= x"2E";
        when x"3853" => data_out<= x"2E";
        when x"3854" => data_out<= x"2E";
        when x"3855" => data_out<= x"00";
        when x"3856" => data_out<= x"49";
        when x"3857" => data_out<= x"6E";
        when x"3858" => data_out<= x"69";
        when x"3859" => data_out<= x"63";
        when x"385A" => data_out<= x"69";
        when x"385B" => data_out<= x"65";
        when x"385C" => data_out<= x"20";
        when x"385D" => data_out<= x"74";
        when x"385E" => data_out<= x"72";
        when x"385F" => data_out<= x"61";
        when x"3860" => data_out<= x"6E";
        when x"3861" => data_out<= x"73";
        when x"3862" => data_out<= x"66";
        when x"3863" => data_out<= x"65";
        when x"3864" => data_out<= x"72";
        when x"3865" => data_out<= x"65";
        when x"3866" => data_out<= x"6E";
        when x"3867" => data_out<= x"63";
        when x"3868" => data_out<= x"69";
        when x"3869" => data_out<= x"61";
        when x"386A" => data_out<= x"2E";
        when x"386B" => data_out<= x"2E";
        when x"386C" => data_out<= x"2E";
        when x"386D" => data_out<= x"00";
        when x"386E" => data_out<= x"45";
        when x"386F" => data_out<= x"6A";
        when x"3870" => data_out<= x"3A";
        when x"3871" => data_out<= x"20";
        when x"3872" => data_out<= x"58";
        when x"3873" => data_out<= x"52";
        when x"3874" => data_out<= x"45";
        when x"3875" => data_out<= x"43";
        when x"3876" => data_out<= x"56";
        when x"3877" => data_out<= x"2C";
        when x"3878" => data_out<= x"20";
        when x"3879" => data_out<= x"58";
        when x"387A" => data_out<= x"52";
        when x"387B" => data_out<= x"45";
        when x"387C" => data_out<= x"43";
        when x"387D" => data_out<= x"56";
        when x"387E" => data_out<= x"20";
        when x"387F" => data_out<= x"31";
        when x"3880" => data_out<= x"30";
        when x"3881" => data_out<= x"30";
        when x"3882" => data_out<= x"30";
        when x"3883" => data_out<= x"0D";
        when x"3884" => data_out<= x"0A";
        when x"3885" => data_out<= x"00";
        when x"3886" => data_out<= x"52";
        when x"3887" => data_out<= x"41";
        when x"3888" => data_out<= x"4D";
        when x"3889" => data_out<= x"20";
        when x"388A" => data_out<= x"70";
        when x"388B" => data_out<= x"72";
        when x"388C" => data_out<= x"6F";
        when x"388D" => data_out<= x"67";
        when x"388E" => data_out<= x"3A";
        when x"388F" => data_out<= x"20";
        when x"3890" => data_out<= x"24";
        when x"3891" => data_out<= x"30";
        when x"3892" => data_out<= x"38";
        when x"3893" => data_out<= x"30";
        when x"3894" => data_out<= x"30";
        when x"3895" => data_out<= x"2D";
        when x"3896" => data_out<= x"24";
        when x"3897" => data_out<= x"33";
        when x"3898" => data_out<= x"44";
        when x"3899" => data_out<= x"46";
        when x"389A" => data_out<= x"46";
        when x"389B" => data_out<= x"0D";
        when x"389C" => data_out<= x"0A";
        when x"389D" => data_out<= x"00";
        when x"389E" => data_out<= x"3D";
        when x"389F" => data_out<= x"3D";
        when x"38A0" => data_out<= x"3D";
        when x"38A1" => data_out<= x"20";
        when x"38A2" => data_out<= x"4D";
        when x"38A3" => data_out<= x"41";
        when x"38A4" => data_out<= x"50";
        when x"38A5" => data_out<= x"41";
        when x"38A6" => data_out<= x"20";
        when x"38A7" => data_out<= x"44";
        when x"38A8" => data_out<= x"45";
        when x"38A9" => data_out<= x"20";
        when x"38AA" => data_out<= x"4D";
        when x"38AB" => data_out<= x"45";
        when x"38AC" => data_out<= x"4D";
        when x"38AD" => data_out<= x"4F";
        when x"38AE" => data_out<= x"52";
        when x"38AF" => data_out<= x"49";
        when x"38B0" => data_out<= x"41";
        when x"38B1" => data_out<= x"20";
        when x"38B2" => data_out<= x"3D";
        when x"38B3" => data_out<= x"3D";
        when x"38B4" => data_out<= x"3D";
        when x"38B5" => data_out<= x"00";
        when x"38B6" => data_out<= x"3D";
        when x"38B7" => data_out<= x"3D";
        when x"38B8" => data_out<= x"3D";
        when x"38B9" => data_out<= x"20";
        when x"38BA" => data_out<= x"4D";
        when x"38BB" => data_out<= x"4F";
        when x"38BC" => data_out<= x"4E";
        when x"38BD" => data_out<= x"49";
        when x"38BE" => data_out<= x"54";
        when x"38BF" => data_out<= x"4F";
        when x"38C0" => data_out<= x"52";
        when x"38C1" => data_out<= x"20";
        when x"38C2" => data_out<= x"36";
        when x"38C3" => data_out<= x"35";
        when x"38C4" => data_out<= x"30";
        when x"38C5" => data_out<= x"32";
        when x"38C6" => data_out<= x"20";
        when x"38C7" => data_out<= x"3D";
        when x"38C8" => data_out<= x"3D";
        when x"38C9" => data_out<= x"3D";
        when x"38CA" => data_out<= x"0D";
        when x"38CB" => data_out<= x"0A";
        when x"38CC" => data_out<= x"00";
        when x"38CD" => data_out<= x"52";
        when x"38CE" => data_out<= x"44";
        when x"38CF" => data_out<= x"20";
        when x"38D0" => data_out<= x"61";
        when x"38D1" => data_out<= x"64";
        when x"38D2" => data_out<= x"64";
        when x"38D3" => data_out<= x"72";
        when x"38D4" => data_out<= x"20";
        when x"38D5" => data_out<= x"20";
        when x"38D6" => data_out<= x"20";
        when x"38D7" => data_out<= x"20";
        when x"38D8" => data_out<= x"4C";
        when x"38D9" => data_out<= x"65";
        when x"38DA" => data_out<= x"65";
        when x"38DB" => data_out<= x"72";
        when x"38DC" => data_out<= x"20";
        when x"38DD" => data_out<= x"62";
        when x"38DE" => data_out<= x"79";
        when x"38DF" => data_out<= x"74";
        when x"38E0" => data_out<= x"65";
        when x"38E1" => data_out<= x"0D";
        when x"38E2" => data_out<= x"0A";
        when x"38E3" => data_out<= x"00";
        when x"38E4" => data_out<= x"45";
        when x"38E5" => data_out<= x"6A";
        when x"38E6" => data_out<= x"3A";
        when x"38E7" => data_out<= x"20";
        when x"38E8" => data_out<= x"52";
        when x"38E9" => data_out<= x"44";
        when x"38EA" => data_out<= x"20";
        when x"38EB" => data_out<= x"30";
        when x"38EC" => data_out<= x"32";
        when x"38ED" => data_out<= x"30";
        when x"38EE" => data_out<= x"30";
        when x"38EF" => data_out<= x"2C";
        when x"38F0" => data_out<= x"20";
        when x"38F1" => data_out<= x"52";
        when x"38F2" => data_out<= x"44";
        when x"38F3" => data_out<= x"20";
        when x"38F4" => data_out<= x"43";
        when x"38F5" => data_out<= x"30";
        when x"38F6" => data_out<= x"30";
        when x"38F7" => data_out<= x"30";
        when x"38F8" => data_out<= x"0D";
        when x"38F9" => data_out<= x"0A";
        when x"38FA" => data_out<= x"00";
        when x"38FB" => data_out<= x"4C";
        when x"38FC" => data_out<= x"69";
        when x"38FD" => data_out<= x"73";
        when x"38FE" => data_out<= x"74";
        when x"38FF" => data_out<= x"6F";
        when x"3900" => data_out<= x"20";
        when x"3901" => data_out<= x"70";
        when x"3902" => data_out<= x"61";
        when x"3903" => data_out<= x"72";
        when x"3904" => data_out<= x"61";
        when x"3905" => data_out<= x"20";
        when x"3906" => data_out<= x"58";
        when x"3907" => data_out<= x"4D";
        when x"3908" => data_out<= x"4F";
        when x"3909" => data_out<= x"44";
        when x"390A" => data_out<= x"45";
        when x"390B" => data_out<= x"4D";
        when x"390C" => data_out<= x"20";
        when x"390D" => data_out<= x"65";
        when x"390E" => data_out<= x"6E";
        when x"390F" => data_out<= x"20";
        when x"3910" => data_out<= x"24";
        when x"3911" => data_out<= x"00";
        when x"3912" => data_out<= x"4C";
        when x"3913" => data_out<= x"65";
        when x"3914" => data_out<= x"6E";
        when x"3915" => data_out<= x"20";
        when x"3916" => data_out<= x"69";
        when x"3917" => data_out<= x"6E";
        when x"3918" => data_out<= x"76";
        when x"3919" => data_out<= x"61";
        when x"391A" => data_out<= x"6C";
        when x"391B" => data_out<= x"69";
        when x"391C" => data_out<= x"64";
        when x"391D" => data_out<= x"6F";
        when x"391E" => data_out<= x"20";
        when x"391F" => data_out<= x"28";
        when x"3920" => data_out<= x"31";
        when x"3921" => data_out<= x"2D";
        when x"3922" => data_out<= x"38";
        when x"3923" => data_out<= x"30";
        when x"3924" => data_out<= x"30";
        when x"3925" => data_out<= x"30";
        when x"3926" => data_out<= x"68";
        when x"3927" => data_out<= x"29";
        when x"3928" => data_out<= x"00";
        when x"3929" => data_out<= x"57";
        when x"392A" => data_out<= x"20";
        when x"392B" => data_out<= x"61";
        when x"392C" => data_out<= x"64";
        when x"392D" => data_out<= x"64";
        when x"392E" => data_out<= x"72";
        when x"392F" => data_out<= x"20";
        when x"3930" => data_out<= x"76";
        when x"3931" => data_out<= x"61";
        when x"3932" => data_out<= x"6C";
        when x"3933" => data_out<= x"20";
        when x"3934" => data_out<= x"45";
        when x"3935" => data_out<= x"73";
        when x"3936" => data_out<= x"63";
        when x"3937" => data_out<= x"72";
        when x"3938" => data_out<= x"69";
        when x"3939" => data_out<= x"62";
        when x"393A" => data_out<= x"69";
        when x"393B" => data_out<= x"72";
        when x"393C" => data_out<= x"0D";
        when x"393D" => data_out<= x"0A";
        when x"393E" => data_out<= x"00";
        when x"393F" => data_out<= x"47";
        when x"3940" => data_out<= x"75";
        when x"3941" => data_out<= x"61";
        when x"3942" => data_out<= x"72";
        when x"3943" => data_out<= x"64";
        when x"3944" => data_out<= x"61";
        when x"3945" => data_out<= x"20";
        when x"3946" => data_out<= x"6D";
        when x"3947" => data_out<= x"65";
        when x"3948" => data_out<= x"6D";
        when x"3949" => data_out<= x"6F";
        when x"394A" => data_out<= x"72";
        when x"394B" => data_out<= x"69";
        when x"394C" => data_out<= x"61";
        when x"394D" => data_out<= x"20";
        when x"394E" => data_out<= x"61";
        when x"394F" => data_out<= x"20";
        when x"3950" => data_out<= x"53";
        when x"3951" => data_out<= x"44";
        when x"3952" => data_out<= x"0D";
        when x"3953" => data_out<= x"0A";
        when x"3954" => data_out<= x"00";
        when x"3955" => data_out<= x"44";
        when x"3956" => data_out<= x"20";
        when x"3957" => data_out<= x"61";
        when x"3958" => data_out<= x"64";
        when x"3959" => data_out<= x"64";
        when x"395A" => data_out<= x"72";
        when x"395B" => data_out<= x"20";
        when x"395C" => data_out<= x"6C";
        when x"395D" => data_out<= x"65";
        when x"395E" => data_out<= x"6E";
        when x"395F" => data_out<= x"20";
        when x"3960" => data_out<= x"44";
        when x"3961" => data_out<= x"75";
        when x"3962" => data_out<= x"6D";
        when x"3963" => data_out<= x"70";
        when x"3964" => data_out<= x"20";
        when x"3965" => data_out<= x"68";
        when x"3966" => data_out<= x"65";
        when x"3967" => data_out<= x"78";
        when x"3968" => data_out<= x"0D";
        when x"3969" => data_out<= x"0A";
        when x"396A" => data_out<= x"00";
        when x"396B" => data_out<= x"52";
        when x"396C" => data_out<= x"44";
        when x"396D" => data_out<= x"20";
        when x"396E" => data_out<= x"61";
        when x"396F" => data_out<= x"64";
        when x"3970" => data_out<= x"64";
        when x"3971" => data_out<= x"72";
        when x"3972" => data_out<= x"20";
        when x"3973" => data_out<= x"2D";
        when x"3974" => data_out<= x"20";
        when x"3975" => data_out<= x"4C";
        when x"3976" => data_out<= x"65";
        when x"3977" => data_out<= x"65";
        when x"3978" => data_out<= x"72";
        when x"3979" => data_out<= x"20";
        when x"397A" => data_out<= x"62";
        when x"397B" => data_out<= x"79";
        when x"397C" => data_out<= x"74";
        when x"397D" => data_out<= x"65";
        when x"397E" => data_out<= x"0D";
        when x"397F" => data_out<= x"0A";
        when x"3980" => data_out<= x"00";
        when x"3981" => data_out<= x"27";
        when x"3982" => data_out<= x"20";
        when x"3983" => data_out<= x"6E";
        when x"3984" => data_out<= x"6F";
        when x"3985" => data_out<= x"20";
        when x"3986" => data_out<= x"65";
        when x"3987" => data_out<= x"78";
        when x"3988" => data_out<= x"69";
        when x"3989" => data_out<= x"73";
        when x"398A" => data_out<= x"74";
        when x"398B" => data_out<= x"65";
        when x"398C" => data_out<= x"2E";
        when x"398D" => data_out<= x"20";
        when x"398E" => data_out<= x"55";
        when x"398F" => data_out<= x"73";
        when x"3990" => data_out<= x"61";
        when x"3991" => data_out<= x"20";
        when x"3992" => data_out<= x"48";
        when x"3993" => data_out<= x"0D";
        when x"3994" => data_out<= x"0A";
        when x"3995" => data_out<= x"00";
        when x"3996" => data_out<= x"53";
        when x"3997" => data_out<= x"41";
        when x"3998" => data_out<= x"56";
        when x"3999" => data_out<= x"45";
        when x"399A" => data_out<= x"20";
        when x"399B" => data_out<= x"66";
        when x"399C" => data_out<= x"69";
        when x"399D" => data_out<= x"6C";
        when x"399E" => data_out<= x"65";
        when x"399F" => data_out<= x"20";
        when x"39A0" => data_out<= x"61";
        when x"39A1" => data_out<= x"64";
        when x"39A2" => data_out<= x"64";
        when x"39A3" => data_out<= x"72";
        when x"39A4" => data_out<= x"20";
        when x"39A5" => data_out<= x"6C";
        when x"39A6" => data_out<= x"65";
        when x"39A7" => data_out<= x"6E";
        when x"39A8" => data_out<= x"0D";
        when x"39A9" => data_out<= x"0A";
        when x"39AA" => data_out<= x"00";
        when x"39AB" => data_out<= x"61";
        when x"39AC" => data_out<= x"64";
        when x"39AD" => data_out<= x"64";
        when x"39AE" => data_out<= x"72";
        when x"39AF" => data_out<= x"20";
        when x"39B0" => data_out<= x"64";
        when x"39B1" => data_out<= x"65";
        when x"39B2" => data_out<= x"66";
        when x"39B3" => data_out<= x"61";
        when x"39B4" => data_out<= x"75";
        when x"39B5" => data_out<= x"6C";
        when x"39B6" => data_out<= x"74";
        when x"39B7" => data_out<= x"3D";
        when x"39B8" => data_out<= x"24";
        when x"39B9" => data_out<= x"30";
        when x"39BA" => data_out<= x"38";
        when x"39BB" => data_out<= x"30";
        when x"39BC" => data_out<= x"30";
        when x"39BD" => data_out<= x"0D";
        when x"39BE" => data_out<= x"0A";
        when x"39BF" => data_out<= x"00";
        when x"39C0" => data_out<= x"4D";
        when x"39C1" => data_out<= x"61";
        when x"39C2" => data_out<= x"78";
        when x"39C3" => data_out<= x"20";
        when x"39C4" => data_out<= x"32";
        when x"39C5" => data_out<= x"35";
        when x"39C6" => data_out<= x"35";
        when x"39C7" => data_out<= x"20";
        when x"39C8" => data_out<= x"28";
        when x"39C9" => data_out<= x"46";
        when x"39CA" => data_out<= x"46";
        when x"39CB" => data_out<= x"29";
        when x"39CC" => data_out<= x"20";
        when x"39CD" => data_out<= x"6C";
        when x"39CE" => data_out<= x"69";
        when x"39CF" => data_out<= x"6E";
        when x"39D0" => data_out<= x"65";
        when x"39D1" => data_out<= x"61";
        when x"39D2" => data_out<= x"73";
        when x"39D3" => data_out<= x"00";
        when x"39D4" => data_out<= x"20";
        when x"39D5" => data_out<= x"28";
        when x"39D6" => data_out<= x"74";
        when x"39D7" => data_out<= x"65";
        when x"39D8" => data_out<= x"72";
        when x"39D9" => data_out<= x"6D";
        when x"39DA" => data_out<= x"69";
        when x"39DB" => data_out<= x"6E";
        when x"39DC" => data_out<= x"61";
        when x"39DD" => data_out<= x"72";
        when x"39DE" => data_out<= x"20";
        when x"39DF" => data_out<= x"63";
        when x"39E0" => data_out<= x"6F";
        when x"39E1" => data_out<= x"6E";
        when x"39E2" => data_out<= x"20";
        when x"39E3" => data_out<= x"27";
        when x"39E4" => data_out<= x"2E";
        when x"39E5" => data_out<= x"27";
        when x"39E6" => data_out<= x"29";
        when x"39E7" => data_out<= x"00";
        when x"39E8" => data_out<= x"52";
        when x"39E9" => data_out<= x"41";
        when x"39EA" => data_out<= x"4D";
        when x"39EB" => data_out<= x"20";
        when x"39EC" => data_out<= x"70";
        when x"39ED" => data_out<= x"61";
        when x"39EE" => data_out<= x"72";
        when x"39EF" => data_out<= x"61";
        when x"39F0" => data_out<= x"20";
        when x"39F1" => data_out<= x"70";
        when x"39F2" => data_out<= x"72";
        when x"39F3" => data_out<= x"6F";
        when x"39F4" => data_out<= x"67";
        when x"39F5" => data_out<= x"72";
        when x"39F6" => data_out<= x"61";
        when x"39F7" => data_out<= x"6D";
        when x"39F8" => data_out<= x"61";
        when x"39F9" => data_out<= x"73";
        when x"39FA" => data_out<= x"3A";
        when x"39FB" => data_out<= x"00";
        when x"39FC" => data_out<= x"4D";
        when x"39FD" => data_out<= x"6F";
        when x"39FE" => data_out<= x"6E";
        when x"39FF" => data_out<= x"74";
        when x"3A00" => data_out<= x"61";
        when x"3A01" => data_out<= x"6E";
        when x"3A02" => data_out<= x"64";
        when x"3A03" => data_out<= x"6F";
        when x"3A04" => data_out<= x"20";
        when x"3A05" => data_out<= x"4D";
        when x"3A06" => data_out<= x"69";
        when x"3A07" => data_out<= x"63";
        when x"3A08" => data_out<= x"72";
        when x"3A09" => data_out<= x"6F";
        when x"3A0A" => data_out<= x"46";
        when x"3A0B" => data_out<= x"53";
        when x"3A0C" => data_out<= x"2E";
        when x"3A0D" => data_out<= x"2E";
        when x"3A0E" => data_out<= x"2E";
        when x"3A0F" => data_out<= x"00";
        when x"3A10" => data_out<= x"45";
        when x"3A11" => data_out<= x"6A";
        when x"3A12" => data_out<= x"3A";
        when x"3A13" => data_out<= x"20";
        when x"3A14" => data_out<= x"44";
        when x"3A15" => data_out<= x"45";
        when x"3A16" => data_out<= x"4C";
        when x"3A17" => data_out<= x"20";
        when x"3A18" => data_out<= x"56";
        when x"3A19" => data_out<= x"49";
        when x"3A1A" => data_out<= x"45";
        when x"3A1B" => data_out<= x"4A";
        when x"3A1C" => data_out<= x"4F";
        when x"3A1D" => data_out<= x"2E";
        when x"3A1E" => data_out<= x"42";
        when x"3A1F" => data_out<= x"49";
        when x"3A20" => data_out<= x"4E";
        when x"3A21" => data_out<= x"0D";
        when x"3A22" => data_out<= x"0A";
        when x"3A23" => data_out<= x"00";
        when x"3A24" => data_out<= x"48";
        when x"3A25" => data_out<= x"2F";
        when x"3A26" => data_out<= x"3F";
        when x"3A27" => data_out<= x"2F";
        when x"3A28" => data_out<= x"51";
        when x"3A29" => data_out<= x"20";
        when x"3A2A" => data_out<= x"41";
        when x"3A2B" => data_out<= x"79";
        when x"3A2C" => data_out<= x"75";
        when x"3A2D" => data_out<= x"64";
        when x"3A2E" => data_out<= x"61";
        when x"3A2F" => data_out<= x"2F";
        when x"3A30" => data_out<= x"53";
        when x"3A31" => data_out<= x"61";
        when x"3A32" => data_out<= x"6C";
        when x"3A33" => data_out<= x"69";
        when x"3A34" => data_out<= x"72";
        when x"3A35" => data_out<= x"0D";
        when x"3A36" => data_out<= x"0A";
        when x"3A37" => data_out<= x"00";
        when x"3A38" => data_out<= x"45";
        when x"3A39" => data_out<= x"6A";
        when x"3A3A" => data_out<= x"3A";
        when x"3A3B" => data_out<= x"20";
        when x"3A3C" => data_out<= x"43";
        when x"3A3D" => data_out<= x"41";
        when x"3A3E" => data_out<= x"54";
        when x"3A3F" => data_out<= x"20";
        when x"3A40" => data_out<= x"50";
        when x"3A41" => data_out<= x"52";
        when x"3A42" => data_out<= x"4F";
        when x"3A43" => data_out<= x"47";
        when x"3A44" => data_out<= x"2E";
        when x"3A45" => data_out<= x"42";
        when x"3A46" => data_out<= x"49";
        when x"3A47" => data_out<= x"4E";
        when x"3A48" => data_out<= x"0D";
        when x"3A49" => data_out<= x"0A";
        when x"3A4A" => data_out<= x"00";
        when x"3A4B" => data_out<= x"4C";
        when x"3A4C" => data_out<= x"4F";
        when x"3A4D" => data_out<= x"41";
        when x"3A4E" => data_out<= x"44";
        when x"3A4F" => data_out<= x"20";
        when x"3A50" => data_out<= x"66";
        when x"3A51" => data_out<= x"69";
        when x"3A52" => data_out<= x"6C";
        when x"3A53" => data_out<= x"65";
        when x"3A54" => data_out<= x"20";
        when x"3A55" => data_out<= x"5B";
        when x"3A56" => data_out<= x"61";
        when x"3A57" => data_out<= x"64";
        when x"3A58" => data_out<= x"64";
        when x"3A59" => data_out<= x"72";
        when x"3A5A" => data_out<= x"5D";
        when x"3A5B" => data_out<= x"0D";
        when x"3A5C" => data_out<= x"0A";
        when x"3A5D" => data_out<= x"00";
        when x"3A5E" => data_out<= x"46";
        when x"3A5F" => data_out<= x"6F";
        when x"3A60" => data_out<= x"72";
        when x"3A61" => data_out<= x"6D";
        when x"3A62" => data_out<= x"61";
        when x"3A63" => data_out<= x"74";
        when x"3A64" => data_out<= x"65";
        when x"3A65" => data_out<= x"61";
        when x"3A66" => data_out<= x"6E";
        when x"3A67" => data_out<= x"64";
        when x"3A68" => data_out<= x"6F";
        when x"3A69" => data_out<= x"20";
        when x"3A6A" => data_out<= x"53";
        when x"3A6B" => data_out<= x"44";
        when x"3A6C" => data_out<= x"2E";
        when x"3A6D" => data_out<= x"2E";
        when x"3A6E" => data_out<= x"2E";
        when x"3A6F" => data_out<= x"00";
        when x"3A70" => data_out<= x"20";
        when x"3A71" => data_out<= x"62";
        when x"3A72" => data_out<= x"79";
        when x"3A73" => data_out<= x"74";
        when x"3A74" => data_out<= x"65";
        when x"3A75" => data_out<= x"73";
        when x"3A76" => data_out<= x"20";
        when x"3A77" => data_out<= x"6D";
        when x"3A78" => data_out<= x"6F";
        when x"3A79" => data_out<= x"73";
        when x"3A7A" => data_out<= x"74";
        when x"3A7B" => data_out<= x"72";
        when x"3A7C" => data_out<= x"61";
        when x"3A7D" => data_out<= x"64";
        when x"3A7E" => data_out<= x"6F";
        when x"3A7F" => data_out<= x"73";
        when x"3A80" => data_out<= x"29";
        when x"3A81" => data_out<= x"00";
        when x"3A82" => data_out<= x"46";
        when x"3A83" => data_out<= x"20";
        when x"3A84" => data_out<= x"61";
        when x"3A85" => data_out<= x"64";
        when x"3A86" => data_out<= x"64";
        when x"3A87" => data_out<= x"72";
        when x"3A88" => data_out<= x"20";
        when x"3A89" => data_out<= x"6C";
        when x"3A8A" => data_out<= x"20";
        when x"3A8B" => data_out<= x"76";
        when x"3A8C" => data_out<= x"20";
        when x"3A8D" => data_out<= x"46";
        when x"3A8E" => data_out<= x"69";
        when x"3A8F" => data_out<= x"6C";
        when x"3A90" => data_out<= x"6C";
        when x"3A91" => data_out<= x"0D";
        when x"3A92" => data_out<= x"0A";
        when x"3A93" => data_out<= x"00";
        when x"3A94" => data_out<= x"4F";
        when x"3A95" => data_out<= x"4B";
        when x"3A96" => data_out<= x"3A";
        when x"3A97" => data_out<= x"20";
        when x"3A98" => data_out<= x"53";
        when x"3A99" => data_out<= x"44";
        when x"3A9A" => data_out<= x"20";
        when x"3A9B" => data_out<= x"66";
        when x"3A9C" => data_out<= x"6F";
        when x"3A9D" => data_out<= x"72";
        when x"3A9E" => data_out<= x"6D";
        when x"3A9F" => data_out<= x"61";
        when x"3AA0" => data_out<= x"74";
        when x"3AA1" => data_out<= x"65";
        when x"3AA2" => data_out<= x"61";
        when x"3AA3" => data_out<= x"64";
        when x"3AA4" => data_out<= x"61";
        when x"3AA5" => data_out<= x"00";
        when x"3AA6" => data_out<= x"20";
        when x"3AA7" => data_out<= x"20";
        when x"3AA8" => data_out<= x"46";
        when x"3AA9" => data_out<= x"6F";
        when x"3AAA" => data_out<= x"72";
        when x"3AAB" => data_out<= x"6D";
        when x"3AAC" => data_out<= x"61";
        when x"3AAD" => data_out<= x"74";
        when x"3AAE" => data_out<= x"65";
        when x"3AAF" => data_out<= x"61";
        when x"3AB0" => data_out<= x"6E";
        when x"3AB1" => data_out<= x"64";
        when x"3AB2" => data_out<= x"6F";
        when x"3AB3" => data_out<= x"2E";
        when x"3AB4" => data_out<= x"2E";
        when x"3AB5" => data_out<= x"2E";
        when x"3AB6" => data_out<= x"00";
        when x"3AB7" => data_out<= x"20";
        when x"3AB8" => data_out<= x"20";
        when x"3AB9" => data_out<= x"53";
        when x"3ABA" => data_out<= x"44";
        when x"3ABB" => data_out<= x"20";
        when x"3ABC" => data_out<= x"4F";
        when x"3ABD" => data_out<= x"4B";
        when x"3ABE" => data_out<= x"2C";
        when x"3ABF" => data_out<= x"20";
        when x"3AC0" => data_out<= x"74";
        when x"3AC1" => data_out<= x"69";
        when x"3AC2" => data_out<= x"70";
        when x"3AC3" => data_out<= x"6F";
        when x"3AC4" => data_out<= x"3A";
        when x"3AC5" => data_out<= x"20";
        when x"3AC6" => data_out<= x"00";
        when x"3AC7" => data_out<= x"4E";
        when x"3AC8" => data_out<= x"6F";
        when x"3AC9" => data_out<= x"20";
        when x"3ACA" => data_out<= x"65";
        when x"3ACB" => data_out<= x"6E";
        when x"3ACC" => data_out<= x"63";
        when x"3ACD" => data_out<= x"6F";
        when x"3ACE" => data_out<= x"6E";
        when x"3ACF" => data_out<= x"74";
        when x"3AD0" => data_out<= x"72";
        when x"3AD1" => data_out<= x"61";
        when x"3AD2" => data_out<= x"64";
        when x"3AD3" => data_out<= x"6F";
        when x"3AD4" => data_out<= x"3A";
        when x"3AD5" => data_out<= x"20";
        when x"3AD6" => data_out<= x"00";
        when x"3AD7" => data_out<= x"45";
        when x"3AD8" => data_out<= x"6A";
        when x"3AD9" => data_out<= x"65";
        when x"3ADA" => data_out<= x"63";
        when x"3ADB" => data_out<= x"75";
        when x"3ADC" => data_out<= x"74";
        when x"3ADD" => data_out<= x"61";
        when x"3ADE" => data_out<= x"6E";
        when x"3ADF" => data_out<= x"64";
        when x"3AE0" => data_out<= x"6F";
        when x"3AE1" => data_out<= x"20";
        when x"3AE2" => data_out<= x"65";
        when x"3AE3" => data_out<= x"6E";
        when x"3AE4" => data_out<= x"20";
        when x"3AE5" => data_out<= x"24";
        when x"3AE6" => data_out<= x"00";
        when x"3AE7" => data_out<= x"20";
        when x"3AE8" => data_out<= x"20";
        when x"3AE9" => data_out<= x"46";
        when x"3AEA" => data_out<= x"53";
        when x"3AEB" => data_out<= x"20";
        when x"3AEC" => data_out<= x"6D";
        when x"3AED" => data_out<= x"6F";
        when x"3AEE" => data_out<= x"6E";
        when x"3AEF" => data_out<= x"74";
        when x"3AF0" => data_out<= x"61";
        when x"3AF1" => data_out<= x"64";
        when x"3AF2" => data_out<= x"6F";
        when x"3AF3" => data_out<= x"20";
        when x"3AF4" => data_out<= x"4F";
        when x"3AF5" => data_out<= x"4B";
        when x"3AF6" => data_out<= x"00";
        when x"3AF7" => data_out<= x"55";
        when x"3AF8" => data_out<= x"73";
        when x"3AF9" => data_out<= x"6F";
        when x"3AFA" => data_out<= x"3A";
        when x"3AFB" => data_out<= x"20";
        when x"3AFC" => data_out<= x"43";
        when x"3AFD" => data_out<= x"41";
        when x"3AFE" => data_out<= x"54";
        when x"3AFF" => data_out<= x"20";
        when x"3B00" => data_out<= x"6E";
        when x"3B01" => data_out<= x"6F";
        when x"3B02" => data_out<= x"6D";
        when x"3B03" => data_out<= x"62";
        when x"3B04" => data_out<= x"72";
        when x"3B05" => data_out<= x"65";
        when x"3B06" => data_out<= x"00";
        when x"3B07" => data_out<= x"55";
        when x"3B08" => data_out<= x"73";
        when x"3B09" => data_out<= x"6F";
        when x"3B0A" => data_out<= x"3A";
        when x"3B0B" => data_out<= x"20";
        when x"3B0C" => data_out<= x"44";
        when x"3B0D" => data_out<= x"45";
        when x"3B0E" => data_out<= x"4C";
        when x"3B0F" => data_out<= x"20";
        when x"3B10" => data_out<= x"6E";
        when x"3B11" => data_out<= x"6F";
        when x"3B12" => data_out<= x"6D";
        when x"3B13" => data_out<= x"62";
        when x"3B14" => data_out<= x"72";
        when x"3B15" => data_out<= x"65";
        when x"3B16" => data_out<= x"00";
        when x"3B17" => data_out<= x"4D";
        when x"3B18" => data_out<= x"6F";
        when x"3B19" => data_out<= x"64";
        when x"3B1A" => data_out<= x"6F";
        when x"3B1B" => data_out<= x"20";
        when x"3B1C" => data_out<= x"63";
        when x"3B1D" => data_out<= x"61";
        when x"3B1E" => data_out<= x"72";
        when x"3B1F" => data_out<= x"67";
        when x"3B20" => data_out<= x"61";
        when x"3B21" => data_out<= x"20";
        when x"3B22" => data_out<= x"65";
        when x"3B23" => data_out<= x"6E";
        when x"3B24" => data_out<= x"20";
        when x"3B25" => data_out<= x"24";
        when x"3B26" => data_out<= x"00";
        when x"3B27" => data_out<= x"20";
        when x"3B28" => data_out<= x"20";
        when x"3B29" => data_out<= x"24";
        when x"3B2A" => data_out<= x"30";
        when x"3B2B" => data_out<= x"38";
        when x"3B2C" => data_out<= x"30";
        when x"3B2D" => data_out<= x"30";
        when x"3B2E" => data_out<= x"2D";
        when x"3B2F" => data_out<= x"24";
        when x"3B30" => data_out<= x"33";
        when x"3B31" => data_out<= x"44";
        when x"3B32" => data_out<= x"46";
        when x"3B33" => data_out<= x"46";
        when x"3B34" => data_out<= x"20";
        when x"3B35" => data_out<= x"28";
        when x"3B36" => data_out<= x"00";
        when x"3B37" => data_out<= x"45";
        when x"3B38" => data_out<= x"72";
        when x"3B39" => data_out<= x"72";
        when x"3B3A" => data_out<= x"6F";
        when x"3B3B" => data_out<= x"72";
        when x"3B3C" => data_out<= x"20";
        when x"3B3D" => data_out<= x"58";
        when x"3B3E" => data_out<= x"4D";
        when x"3B3F" => data_out<= x"4F";
        when x"3B40" => data_out<= x"44";
        when x"3B41" => data_out<= x"45";
        when x"3B42" => data_out<= x"4D";
        when x"3B43" => data_out<= x"3A";
        when x"3B44" => data_out<= x"20";
        when x"3B45" => data_out<= x"00";
        when x"3B46" => data_out<= x"53";
        when x"3B47" => data_out<= x"44";
        when x"3B48" => data_out<= x"20";
        when x"3B49" => data_out<= x"6E";
        when x"3B4A" => data_out<= x"6F";
        when x"3B4B" => data_out<= x"20";
        when x"3B4C" => data_out<= x"6D";
        when x"3B4D" => data_out<= x"6F";
        when x"3B4E" => data_out<= x"6E";
        when x"3B4F" => data_out<= x"74";
        when x"3B50" => data_out<= x"61";
        when x"3B51" => data_out<= x"64";
        when x"3B52" => data_out<= x"61";
        when x"3B53" => data_out<= x"00";
        when x"3B54" => data_out<= x"4E";
        when x"3B55" => data_out<= x"6F";
        when x"3B56" => data_out<= x"20";
        when x"3B57" => data_out<= x"65";
        when x"3B58" => data_out<= x"6E";
        when x"3B59" => data_out<= x"63";
        when x"3B5A" => data_out<= x"6F";
        when x"3B5B" => data_out<= x"6E";
        when x"3B5C" => data_out<= x"74";
        when x"3B5D" => data_out<= x"72";
        when x"3B5E" => data_out<= x"61";
        when x"3B5F" => data_out<= x"64";
        when x"3B60" => data_out<= x"6F";
        when x"3B61" => data_out<= x"00";
        when x"3B62" => data_out<= x"45";
        when x"3B63" => data_out<= x"72";
        when x"3B64" => data_out<= x"72";
        when x"3B65" => data_out<= x"6F";
        when x"3B66" => data_out<= x"72";
        when x"3B67" => data_out<= x"20";
        when x"3B68" => data_out<= x"63";
        when x"3B69" => data_out<= x"72";
        when x"3B6A" => data_out<= x"65";
        when x"3B6B" => data_out<= x"61";
        when x"3B6C" => data_out<= x"72";
        when x"3B6D" => data_out<= x"3A";
        when x"3B6E" => data_out<= x"20";
        when x"3B6F" => data_out<= x"00";
        when x"3B70" => data_out<= x"2F";
        when x"3B71" => data_out<= x"31";
        when x"3B72" => data_out<= x"36";
        when x"3B73" => data_out<= x"20";
        when x"3B74" => data_out<= x"61";
        when x"3B75" => data_out<= x"72";
        when x"3B76" => data_out<= x"63";
        when x"3B77" => data_out<= x"68";
        when x"3B78" => data_out<= x"69";
        when x"3B79" => data_out<= x"76";
        when x"3B7A" => data_out<= x"6F";
        when x"3B7B" => data_out<= x"73";
        when x"3B7C" => data_out<= x"00";
        when x"3B7D" => data_out<= x"2D";
        when x"3B7E" => data_out<= x"2D";
        when x"3B7F" => data_out<= x"2D";
        when x"3B80" => data_out<= x"20";
        when x"3B81" => data_out<= x"53";
        when x"3B82" => data_out<= x"44";
        when x"3B83" => data_out<= x"20";
        when x"3B84" => data_out<= x"2D";
        when x"3B85" => data_out<= x"2D";
        when x"3B86" => data_out<= x"2D";
        when x"3B87" => data_out<= x"0D";
        when x"3B88" => data_out<= x"0A";
        when x"3B89" => data_out<= x"00";
        when x"3B8A" => data_out<= x"20";
        when x"3B8B" => data_out<= x"62";
        when x"3B8C" => data_out<= x"79";
        when x"3B8D" => data_out<= x"74";
        when x"3B8E" => data_out<= x"65";
        when x"3B8F" => data_out<= x"73";
        when x"3B90" => data_out<= x"29";
        when x"3B91" => data_out<= x"20";
        when x"3B92" => data_out<= x"2D";
        when x"3B93" => data_out<= x"3E";
        when x"3B94" => data_out<= x"20";
        when x"3B95" => data_out<= x"24";
        when x"3B96" => data_out<= x"00";
        when x"3B97" => data_out<= x"52";
        when x"3B98" => data_out<= x"65";
        when x"3B99" => data_out<= x"74";
        when x"3B9A" => data_out<= x"6F";
        when x"3B9B" => data_out<= x"72";
        when x"3B9C" => data_out<= x"6E";
        when x"3B9D" => data_out<= x"6F";
        when x"3B9E" => data_out<= x"20";
        when x"3B9F" => data_out<= x"64";
        when x"3BA0" => data_out<= x"65";
        when x"3BA1" => data_out<= x"20";
        when x"3BA2" => data_out<= x"24";
        when x"3BA3" => data_out<= x"00";
        when x"3BA4" => data_out<= x"20";
        when x"3BA5" => data_out<= x"20";
        when x"3BA6" => data_out<= x"45";
        when x"3BA7" => data_out<= x"72";
        when x"3BA8" => data_out<= x"72";
        when x"3BA9" => data_out<= x"6F";
        when x"3BAA" => data_out<= x"72";
        when x"3BAB" => data_out<= x"20";
        when x"3BAC" => data_out<= x"53";
        when x"3BAD" => data_out<= x"44";
        when x"3BAE" => data_out<= x"3A";
        when x"3BAF" => data_out<= x"20";
        when x"3BB0" => data_out<= x"00";
        when x"3BB1" => data_out<= x"20";
        when x"3BB2" => data_out<= x"20";
        when x"3BB3" => data_out<= x"45";
        when x"3BB4" => data_out<= x"72";
        when x"3BB5" => data_out<= x"72";
        when x"3BB6" => data_out<= x"6F";
        when x"3BB7" => data_out<= x"72";
        when x"3BB8" => data_out<= x"20";
        when x"3BB9" => data_out<= x"46";
        when x"3BBA" => data_out<= x"53";
        when x"3BBB" => data_out<= x"3A";
        when x"3BBC" => data_out<= x"20";
        when x"3BBD" => data_out<= x"00";
        when x"3BBE" => data_out<= x"47";
        when x"3BBF" => data_out<= x"75";
        when x"3BC0" => data_out<= x"61";
        when x"3BC1" => data_out<= x"72";
        when x"3BC2" => data_out<= x"64";
        when x"3BC3" => data_out<= x"61";
        when x"3BC4" => data_out<= x"6E";
        when x"3BC5" => data_out<= x"64";
        when x"3BC6" => data_out<= x"6F";
        when x"3BC7" => data_out<= x"20";
        when x"3BC8" => data_out<= x"24";
        when x"3BC9" => data_out<= x"00";
        when x"3BCA" => data_out<= x"20";
        when x"3BCB" => data_out<= x"62";
        when x"3BCC" => data_out<= x"79";
        when x"3BCD" => data_out<= x"74";
        when x"3BCE" => data_out<= x"65";
        when x"3BCF" => data_out<= x"73";
        when x"3BD0" => data_out<= x"20";
        when x"3BD1" => data_out<= x"65";
        when x"3BD2" => data_out<= x"6E";
        when x"3BD3" => data_out<= x"20";
        when x"3BD4" => data_out<= x"24";
        when x"3BD5" => data_out<= x"00";
        when x"3BD6" => data_out<= x"45";
        when x"3BD7" => data_out<= x"6C";
        when x"3BD8" => data_out<= x"69";
        when x"3BD9" => data_out<= x"6D";
        when x"3BDA" => data_out<= x"69";
        when x"3BDB" => data_out<= x"6E";
        when x"3BDC" => data_out<= x"61";
        when x"3BDD" => data_out<= x"64";
        when x"3BDE" => data_out<= x"6F";
        when x"3BDF" => data_out<= x"3A";
        when x"3BE0" => data_out<= x"20";
        when x"3BE1" => data_out<= x"00";
        when x"3BE2" => data_out<= x"43";
        when x"3BE3" => data_out<= x"61";
        when x"3BE4" => data_out<= x"72";
        when x"3BE5" => data_out<= x"67";
        when x"3BE6" => data_out<= x"61";
        when x"3BE7" => data_out<= x"64";
        when x"3BE8" => data_out<= x"6F";
        when x"3BE9" => data_out<= x"73";
        when x"3BEA" => data_out<= x"20";
        when x"3BEB" => data_out<= x"00";
        when x"3BEC" => data_out<= x"43";
        when x"3BED" => data_out<= x"61";
        when x"3BEE" => data_out<= x"72";
        when x"3BEF" => data_out<= x"67";
        when x"3BF0" => data_out<= x"61";
        when x"3BF1" => data_out<= x"6E";
        when x"3BF2" => data_out<= x"64";
        when x"3BF3" => data_out<= x"6F";
        when x"3BF4" => data_out<= x"20";
        when x"3BF5" => data_out<= x"00";
        when x"3BF6" => data_out<= x"20";
        when x"3BF7" => data_out<= x"20";
        when x"3BF8" => data_out<= x"28";
        when x"3BF9" => data_out<= x"76";
        when x"3BFA" => data_out<= x"61";
        when x"3BFB" => data_out<= x"63";
        when x"3BFC" => data_out<= x"69";
        when x"3BFD" => data_out<= x"6F";
        when x"3BFE" => data_out<= x"29";
        when x"3BFF" => data_out<= x"00";
        when x"3C00" => data_out<= x"41";
        when x"3C01" => data_out<= x"72";
        when x"3C02" => data_out<= x"63";
        when x"3C03" => data_out<= x"68";
        when x"3C04" => data_out<= x"69";
        when x"3C05" => data_out<= x"76";
        when x"3C06" => data_out<= x"6F";
        when x"3C07" => data_out<= x"73";
        when x"3C08" => data_out<= x"3A";
        when x"3C09" => data_out<= x"00";
        when x"3C0A" => data_out<= x"53";
        when x"3C0B" => data_out<= x"44";
        when x"3C0C" => data_out<= x"46";
        when x"3C0D" => data_out<= x"4F";
        when x"3C0E" => data_out<= x"52";
        when x"3C0F" => data_out<= x"4D";
        when x"3C10" => data_out<= x"41";
        when x"3C11" => data_out<= x"54";
        when x"3C12" => data_out<= x"00";
        when x"3C13" => data_out<= x"46";
        when x"3C14" => data_out<= x"69";
        when x"3C15" => data_out<= x"6C";
        when x"3C16" => data_out<= x"6C";
        when x"3C17" => data_out<= x"65";
        when x"3C18" => data_out<= x"64";
        when x"3C19" => data_out<= x"20";
        when x"3C1A" => data_out<= x"24";
        when x"3C1B" => data_out<= x"00";
        when x"3C1C" => data_out<= x"20";
        when x"3C1D" => data_out<= x"62";
        when x"3C1E" => data_out<= x"79";
        when x"3C1F" => data_out<= x"74";
        when x"3C20" => data_out<= x"65";
        when x"3C21" => data_out<= x"73";
        when x"3C22" => data_out<= x"29";
        when x"3C23" => data_out<= x"00";
        when x"3C24" => data_out<= x"54";
        when x"3C25" => data_out<= x"6F";
        when x"3C26" => data_out<= x"74";
        when x"3C27" => data_out<= x"61";
        when x"3C28" => data_out<= x"6C";
        when x"3C29" => data_out<= x"3A";
        when x"3C2A" => data_out<= x"20";
        when x"3C2B" => data_out<= x"00";
        when x"3C2C" => data_out<= x"45";
        when x"3C2D" => data_out<= x"72";
        when x"3C2E" => data_out<= x"72";
        when x"3C2F" => data_out<= x"6F";
        when x"3C30" => data_out<= x"72";
        when x"3C31" => data_out<= x"3A";
        when x"3C32" => data_out<= x"20";
        when x"3C33" => data_out<= x"00";
        when x"3C34" => data_out<= x"20";
        when x"3C35" => data_out<= x"62";
        when x"3C36" => data_out<= x"79";
        when x"3C37" => data_out<= x"74";
        when x"3C38" => data_out<= x"65";
        when x"3C39" => data_out<= x"73";
        when x"3C3A" => data_out<= x"00";
        when x"3C3B" => data_out<= x"20";
        when x"3C3C" => data_out<= x"5B";
        when x"3C3D" => data_out<= x"45";
        when x"3C3E" => data_out<= x"53";
        when x"3C3F" => data_out<= x"43";
        when x"3C40" => data_out<= x"5D";
        when x"3C41" => data_out<= x"00";
        when x"3C42" => data_out<= x"20";
        when x"3C43" => data_out<= x"63";
        when x"3C44" => data_out<= x"6F";
        when x"3C45" => data_out<= x"6E";
        when x"3C46" => data_out<= x"20";
        when x"3C47" => data_out<= x"24";
        when x"3C48" => data_out<= x"00";
        when x"3C49" => data_out<= x"43";
        when x"3C4A" => data_out<= x"6D";
        when x"3C4B" => data_out<= x"64";
        when x"3C4C" => data_out<= x"20";
        when x"3C4D" => data_out<= x"27";
        when x"3C4E" => data_out<= x"00";
        when x"3C4F" => data_out<= x"4C";
        when x"3C50" => data_out<= x"44";
        when x"3C51" => data_out<= x"41";
        when x"3C52" => data_out<= x"7A";
        when x"3C53" => data_out<= x"70";
        when x"3C54" => data_out<= x"00";
        when x"3C55" => data_out<= x"20";
        when x"3C56" => data_out<= x"3C";
        when x"3C57" => data_out<= x"2D";
        when x"3C58" => data_out<= x"20";
        when x"3C59" => data_out<= x"24";
        when x"3C5A" => data_out<= x"00";
        when x"3C5B" => data_out<= x"4C";
        when x"3C5C" => data_out<= x"44";
        when x"3C5D" => data_out<= x"41";
        when x"3C5E" => data_out<= x"61";
        when x"3C5F" => data_out<= x"62";
        when x"3C60" => data_out<= x"00";
        when x"3C61" => data_out<= x"58";
        when x"3C62" => data_out<= x"52";
        when x"3C63" => data_out<= x"45";
        when x"3C64" => data_out<= x"43";
        when x"3C65" => data_out<= x"56";
        when x"3C66" => data_out<= x"00";
        when x"3C67" => data_out<= x"4A";
        when x"3C68" => data_out<= x"4D";
        when x"3C69" => data_out<= x"50";
        when x"3C6A" => data_out<= x"28";
        when x"3C6B" => data_out<= x"29";
        when x"3C6C" => data_out<= x"00";
        when x"3C6D" => data_out<= x"53";
        when x"3C6E" => data_out<= x"54";
        when x"3C6F" => data_out<= x"41";
        when x"3C70" => data_out<= x"7A";
        when x"3C71" => data_out<= x"70";
        when x"3C72" => data_out<= x"00";
        when x"3C73" => data_out<= x"53";
        when x"3C74" => data_out<= x"54";
        when x"3C75" => data_out<= x"41";
        when x"3C76" => data_out<= x"61";
        when x"3C77" => data_out<= x"62";
        when x"3C78" => data_out<= x"00";
        when x"3C79" => data_out<= x"53";
        when x"3C7A" => data_out<= x"54";
        when x"3C7B" => data_out<= x"58";
        when x"3C7C" => data_out<= x"7A";
        when x"3C7D" => data_out<= x"70";
        when x"3C7E" => data_out<= x"00";
        when x"3C7F" => data_out<= x"45";
        when x"3C80" => data_out<= x"52";
        when x"3C81" => data_out<= x"52";
        when x"3C82" => data_out<= x"3A";
        when x"3C83" => data_out<= x"20";
        when x"3C84" => data_out<= x"00";
        when x"3C85" => data_out<= x"53";
        when x"3C86" => data_out<= x"54";
        when x"3C87" => data_out<= x"59";
        when x"3C88" => data_out<= x"7A";
        when x"3C89" => data_out<= x"70";
        when x"3C8A" => data_out<= x"00";
        when x"3C8B" => data_out<= x"20";
        when x"3C8C" => data_out<= x"2D";
        when x"3C8D" => data_out<= x"3E";
        when x"3C8E" => data_out<= x"20";
        when x"3C8F" => data_out<= x"00";
        when x"3C90" => data_out<= x"4C";
        when x"3C91" => data_out<= x"44";
        when x"3C92" => data_out<= x"41";
        when x"3C93" => data_out<= x"23";
        when x"3C94" => data_out<= x"00";
        when x"3C95" => data_out<= x"4C";
        when x"3C96" => data_out<= x"4F";
        when x"3C97" => data_out<= x"41";
        when x"3C98" => data_out<= x"44";
        when x"3C99" => data_out<= x"00";
        when x"3C9A" => data_out<= x"53";
        when x"3C9B" => data_out<= x"41";
        when x"3C9C" => data_out<= x"56";
        when x"3C9D" => data_out<= x"45";
        when x"3C9E" => data_out<= x"00";
        when x"3C9F" => data_out<= x"20";
        when x"3CA0" => data_out<= x"3D";
        when x"3CA1" => data_out<= x"20";
        when x"3CA2" => data_out<= x"24";
        when x"3CA3" => data_out<= x"00";
        when x"3CA4" => data_out<= x"4F";
        when x"3CA5" => data_out<= x"4B";
        when x"3CA6" => data_out<= x"3A";
        when x"3CA7" => data_out<= x"20";
        when x"3CA8" => data_out<= x"00";
        when x"3CA9" => data_out<= x"41";
        when x"3CAA" => data_out<= x"44";
        when x"3CAB" => data_out<= x"43";
        when x"3CAC" => data_out<= x"23";
        when x"3CAD" => data_out<= x"00";
        when x"3CAE" => data_out<= x"45";
        when x"3CAF" => data_out<= x"4F";
        when x"3CB0" => data_out<= x"52";
        when x"3CB1" => data_out<= x"23";
        when x"3CB2" => data_out<= x"00";
        when x"3CB3" => data_out<= x"4F";
        when x"3CB4" => data_out<= x"52";
        when x"3CB5" => data_out<= x"41";
        when x"3CB6" => data_out<= x"23";
        when x"3CB7" => data_out<= x"00";
        when x"3CB8" => data_out<= x"3D";
        when x"3CB9" => data_out<= x"3D";
        when x"3CBA" => data_out<= x"3D";
        when x"3CBB" => data_out<= x"20";
        when x"3CBC" => data_out<= x"00";
        when x"3CBD" => data_out<= x"4C";
        when x"3CBE" => data_out<= x"44";
        when x"3CBF" => data_out<= x"58";
        when x"3CC0" => data_out<= x"23";
        when x"3CC1" => data_out<= x"00";
        when x"3CC2" => data_out<= x"4C";
        when x"3CC3" => data_out<= x"44";
        when x"3CC4" => data_out<= x"59";
        when x"3CC5" => data_out<= x"23";
        when x"3CC6" => data_out<= x"00";
        when x"3CC7" => data_out<= x"2E";
        when x"3CC8" => data_out<= x"2E";
        when x"3CC9" => data_out<= x"2E";
        when x"3CCA" => data_out<= x"28";
        when x"3CCB" => data_out<= x"00";
        when x"3CCC" => data_out<= x"41";
        when x"3CCD" => data_out<= x"4E";
        when x"3CCE" => data_out<= x"44";
        when x"3CCF" => data_out<= x"23";
        when x"3CD0" => data_out<= x"00";
        when x"3CD1" => data_out<= x"43";
        when x"3CD2" => data_out<= x"50";
        when x"3CD3" => data_out<= x"59";
        when x"3CD4" => data_out<= x"23";
        when x"3CD5" => data_out<= x"00";
        when x"3CD6" => data_out<= x"43";
        when x"3CD7" => data_out<= x"50";
        when x"3CD8" => data_out<= x"58";
        when x"3CD9" => data_out<= x"23";
        when x"3CDA" => data_out<= x"00";
        when x"3CDB" => data_out<= x"43";
        when x"3CDC" => data_out<= x"4D";
        when x"3CDD" => data_out<= x"50";
        when x"3CDE" => data_out<= x"23";
        when x"3CDF" => data_out<= x"00";
        when x"3CE0" => data_out<= x"53";
        when x"3CE1" => data_out<= x"42";
        when x"3CE2" => data_out<= x"43";
        when x"3CE3" => data_out<= x"23";
        when x"3CE4" => data_out<= x"00";
        when x"3CE5" => data_out<= x"49";
        when x"3CE6" => data_out<= x"4E";
        when x"3CE7" => data_out<= x"59";
        when x"3CE8" => data_out<= x"00";
        when x"3CE9" => data_out<= x"49";
        when x"3CEA" => data_out<= x"4E";
        when x"3CEB" => data_out<= x"58";
        when x"3CEC" => data_out<= x"00";
        when x"3CED" => data_out<= x"44";
        when x"3CEE" => data_out<= x"45";
        when x"3CEF" => data_out<= x"59";
        when x"3CF0" => data_out<= x"00";
        when x"3CF1" => data_out<= x"43";
        when x"3CF2" => data_out<= x"4C";
        when x"3CF3" => data_out<= x"43";
        when x"3CF4" => data_out<= x"00";
        when x"3CF5" => data_out<= x"53";
        when x"3CF6" => data_out<= x"45";
        when x"3CF7" => data_out<= x"43";
        when x"3CF8" => data_out<= x"00";
        when x"3CF9" => data_out<= x"43";
        when x"3CFA" => data_out<= x"4C";
        when x"3CFB" => data_out<= x"44";
        when x"3CFC" => data_out<= x"00";
        when x"3CFD" => data_out<= x"53";
        when x"3CFE" => data_out<= x"45";
        when x"3CFF" => data_out<= x"44";
        when x"3D00" => data_out<= x"00";
        when x"3D01" => data_out<= x"20";
        when x"3D02" => data_out<= x"20";
        when x"3D03" => data_out<= x"20";
        when x"3D04" => data_out<= x"00";
        when x"3D05" => data_out<= x"42";
        when x"3D06" => data_out<= x"4E";
        when x"3D07" => data_out<= x"45";
        when x"3D08" => data_out<= x"00";
        when x"3D09" => data_out<= x"42";
        when x"3D0A" => data_out<= x"45";
        when x"3D0B" => data_out<= x"51";
        when x"3D0C" => data_out<= x"00";
        when x"3D0D" => data_out<= x"42";
        when x"3D0E" => data_out<= x"50";
        when x"3D0F" => data_out<= x"4C";
        when x"3D10" => data_out<= x"00";
        when x"3D11" => data_out<= x"44";
        when x"3D12" => data_out<= x"45";
        when x"3D13" => data_out<= x"4C";
        when x"3D14" => data_out<= x"00";
        when x"3D15" => data_out<= x"43";
        when x"3D16" => data_out<= x"4C";
        when x"3D17" => data_out<= x"49";
        when x"3D18" => data_out<= x"00";
        when x"3D19" => data_out<= x"4A";
        when x"3D1A" => data_out<= x"4D";
        when x"3D1B" => data_out<= x"50";
        when x"3D1C" => data_out<= x"00";
        when x"3D1D" => data_out<= x"52";
        when x"3D1E" => data_out<= x"54";
        when x"3D1F" => data_out<= x"53";
        when x"3D20" => data_out<= x"00";
        when x"3D21" => data_out<= x"52";
        when x"3D22" => data_out<= x"54";
        when x"3D23" => data_out<= x"49";
        when x"3D24" => data_out<= x"00";
        when x"3D25" => data_out<= x"4A";
        when x"3D26" => data_out<= x"53";
        when x"3D27" => data_out<= x"52";
        when x"3D28" => data_out<= x"00";
        when x"3D29" => data_out<= x"42";
        when x"3D2A" => data_out<= x"52";
        when x"3D2B" => data_out<= x"4B";
        when x"3D2C" => data_out<= x"00";
        when x"3D2D" => data_out<= x"42";
        when x"3D2E" => data_out<= x"4D";
        when x"3D2F" => data_out<= x"49";
        when x"3D30" => data_out<= x"00";
        when x"3D31" => data_out<= x"42";
        when x"3D32" => data_out<= x"43";
        when x"3D33" => data_out<= x"43";
        when x"3D34" => data_out<= x"00";
        when x"3D35" => data_out<= x"53";
        when x"3D36" => data_out<= x"45";
        when x"3D37" => data_out<= x"49";
        when x"3D38" => data_out<= x"00";
        when x"3D39" => data_out<= x"43";
        when x"3D3A" => data_out<= x"41";
        when x"3D3B" => data_out<= x"54";
        when x"3D3C" => data_out<= x"00";
        when x"3D3D" => data_out<= x"4E";
        when x"3D3E" => data_out<= x"4F";
        when x"3D3F" => data_out<= x"50";
        when x"3D40" => data_out<= x"00";
        when x"3D41" => data_out<= x"54";
        when x"3D42" => data_out<= x"41";
        when x"3D43" => data_out<= x"58";
        when x"3D44" => data_out<= x"00";
        when x"3D45" => data_out<= x"42";
        when x"3D46" => data_out<= x"43";
        when x"3D47" => data_out<= x"53";
        when x"3D48" => data_out<= x"00";
        when x"3D49" => data_out<= x"54";
        when x"3D4A" => data_out<= x"41";
        when x"3D4B" => data_out<= x"59";
        when x"3D4C" => data_out<= x"00";
        when x"3D4D" => data_out<= x"54";
        when x"3D4E" => data_out<= x"58";
        when x"3D4F" => data_out<= x"41";
        when x"3D50" => data_out<= x"00";
        when x"3D51" => data_out<= x"54";
        when x"3D52" => data_out<= x"59";
        when x"3D53" => data_out<= x"41";
        when x"3D54" => data_out<= x"00";
        when x"3D55" => data_out<= x"42";
        when x"3D56" => data_out<= x"56";
        when x"3D57" => data_out<= x"43";
        when x"3D58" => data_out<= x"00";
        when x"3D59" => data_out<= x"42";
        when x"3D5A" => data_out<= x"56";
        when x"3D5B" => data_out<= x"53";
        when x"3D5C" => data_out<= x"00";
        when x"3D5D" => data_out<= x"54";
        when x"3D5E" => data_out<= x"58";
        when x"3D5F" => data_out<= x"53";
        when x"3D60" => data_out<= x"00";
        when x"3D61" => data_out<= x"3F";
        when x"3D62" => data_out<= x"3F";
        when x"3D63" => data_out<= x"3F";
        when x"3D64" => data_out<= x"00";
        when x"3D65" => data_out<= x"54";
        when x"3D66" => data_out<= x"53";
        when x"3D67" => data_out<= x"58";
        when x"3D68" => data_out<= x"00";
        when x"3D69" => data_out<= x"50";
        when x"3D6A" => data_out<= x"48";
        when x"3D6B" => data_out<= x"41";
        when x"3D6C" => data_out<= x"00";
        when x"3D6D" => data_out<= x"50";
        when x"3D6E" => data_out<= x"4C";
        when x"3D6F" => data_out<= x"41";
        when x"3D70" => data_out<= x"00";
        when x"3D71" => data_out<= x"50";
        when x"3D72" => data_out<= x"48";
        when x"3D73" => data_out<= x"50";
        when x"3D74" => data_out<= x"00";
        when x"3D75" => data_out<= x"50";
        when x"3D76" => data_out<= x"4C";
        when x"3D77" => data_out<= x"50";
        when x"3D78" => data_out<= x"00";
        when x"3D79" => data_out<= x"44";
        when x"3D7A" => data_out<= x"45";
        when x"3D7B" => data_out<= x"58";
        when x"3D7C" => data_out<= x"00";
        when x"3D7D" => data_out<= x"2D";
        when x"3D7E" => data_out<= x"24";
        when x"3D7F" => data_out<= x"00";
        when x"3D80" => data_out<= x"4C";
        when x"3D81" => data_out<= x"53";
        when x"3D82" => data_out<= x"00";
        when x"3D83" => data_out<= x"00";
        when x"3D84" => data_out<= x"00";
        when x"3D85" => data_out<= x"00";
        when x"3D86" => data_out<= x"02";
        when x"3D87" => data_out<= x"00";
        when x"3D88" => data_out<= x"00";
        when x"3D89" => data_out<= x"00";
        when x"3D8A" => data_out<= x"00";
        when x"3D8B" => data_out<= x"EA";
        when x"3D8C" => data_out<= x"EA";
        when x"3D8D" => data_out<= x"EA";
        when x"3D8E" => data_out<= x"EA";
        when x"3D8F" => data_out<= x"EA";
        when x"3D90" => data_out<= x"EA";
        when x"3D91" => data_out<= x"EA";
        when x"3D92" => data_out<= x"EA";
        when x"3D93" => data_out<= x"EA";
        when x"3D94" => data_out<= x"EA";
        when x"3D95" => data_out<= x"EA";
        when x"3D96" => data_out<= x"EA";
        when x"3D97" => data_out<= x"EA";
        when x"3D98" => data_out<= x"EA";
        when x"3D99" => data_out<= x"EA";
        when x"3D9A" => data_out<= x"EA";
        when x"3D9B" => data_out<= x"EA";
        when x"3D9C" => data_out<= x"EA";
        when x"3D9D" => data_out<= x"EA";
        when x"3D9E" => data_out<= x"EA";
        when x"3D9F" => data_out<= x"EA";
        when x"3DA0" => data_out<= x"EA";
        when x"3DA1" => data_out<= x"EA";
        when x"3DA2" => data_out<= x"EA";
        when x"3DA3" => data_out<= x"EA";
        when x"3DA4" => data_out<= x"EA";
        when x"3DA5" => data_out<= x"EA";
        when x"3DA6" => data_out<= x"EA";
        when x"3DA7" => data_out<= x"EA";
        when x"3DA8" => data_out<= x"EA";
        when x"3DA9" => data_out<= x"EA";
        when x"3DAA" => data_out<= x"EA";
        when x"3DAB" => data_out<= x"EA";
        when x"3DAC" => data_out<= x"EA";
        when x"3DAD" => data_out<= x"EA";
        when x"3DAE" => data_out<= x"EA";
        when x"3DAF" => data_out<= x"EA";
        when x"3DB0" => data_out<= x"EA";
        when x"3DB1" => data_out<= x"EA";
        when x"3DB2" => data_out<= x"EA";
        when x"3DB3" => data_out<= x"EA";
        when x"3DB4" => data_out<= x"EA";
        when x"3DB5" => data_out<= x"EA";
        when x"3DB6" => data_out<= x"EA";
        when x"3DB7" => data_out<= x"EA";
        when x"3DB8" => data_out<= x"EA";
        when x"3DB9" => data_out<= x"EA";
        when x"3DBA" => data_out<= x"EA";
        when x"3DBB" => data_out<= x"EA";
        when x"3DBC" => data_out<= x"EA";
        when x"3DBD" => data_out<= x"EA";
        when x"3DBE" => data_out<= x"EA";
        when x"3DBF" => data_out<= x"EA";
        when x"3DC0" => data_out<= x"EA";
        when x"3DC1" => data_out<= x"EA";
        when x"3DC2" => data_out<= x"EA";
        when x"3DC3" => data_out<= x"EA";
        when x"3DC4" => data_out<= x"EA";
        when x"3DC5" => data_out<= x"EA";
        when x"3DC6" => data_out<= x"EA";
        when x"3DC7" => data_out<= x"EA";
        when x"3DC8" => data_out<= x"EA";
        when x"3DC9" => data_out<= x"EA";
        when x"3DCA" => data_out<= x"EA";
        when x"3DCB" => data_out<= x"EA";
        when x"3DCC" => data_out<= x"EA";
        when x"3DCD" => data_out<= x"EA";
        when x"3DCE" => data_out<= x"EA";
        when x"3DCF" => data_out<= x"EA";
        when x"3DD0" => data_out<= x"EA";
        when x"3DD1" => data_out<= x"EA";
        when x"3DD2" => data_out<= x"EA";
        when x"3DD3" => data_out<= x"EA";
        when x"3DD4" => data_out<= x"EA";
        when x"3DD5" => data_out<= x"EA";
        when x"3DD6" => data_out<= x"EA";
        when x"3DD7" => data_out<= x"EA";
        when x"3DD8" => data_out<= x"EA";
        when x"3DD9" => data_out<= x"EA";
        when x"3DDA" => data_out<= x"EA";
        when x"3DDB" => data_out<= x"EA";
        when x"3DDC" => data_out<= x"EA";
        when x"3DDD" => data_out<= x"EA";
        when x"3DDE" => data_out<= x"EA";
        when x"3DDF" => data_out<= x"EA";
        when x"3DE0" => data_out<= x"EA";
        when x"3DE1" => data_out<= x"EA";
        when x"3DE2" => data_out<= x"EA";
        when x"3DE3" => data_out<= x"EA";
        when x"3DE4" => data_out<= x"EA";
        when x"3DE5" => data_out<= x"EA";
        when x"3DE6" => data_out<= x"EA";
        when x"3DE7" => data_out<= x"EA";
        when x"3DE8" => data_out<= x"EA";
        when x"3DE9" => data_out<= x"EA";
        when x"3DEA" => data_out<= x"EA";
        when x"3DEB" => data_out<= x"EA";
        when x"3DEC" => data_out<= x"EA";
        when x"3DED" => data_out<= x"EA";
        when x"3DEE" => data_out<= x"EA";
        when x"3DEF" => data_out<= x"EA";
        when x"3DF0" => data_out<= x"EA";
        when x"3DF1" => data_out<= x"EA";
        when x"3DF2" => data_out<= x"EA";
        when x"3DF3" => data_out<= x"EA";
        when x"3DF4" => data_out<= x"EA";
        when x"3DF5" => data_out<= x"EA";
        when x"3DF6" => data_out<= x"EA";
        when x"3DF7" => data_out<= x"EA";
        when x"3DF8" => data_out<= x"EA";
        when x"3DF9" => data_out<= x"EA";
        when x"3DFA" => data_out<= x"EA";
        when x"3DFB" => data_out<= x"EA";
        when x"3DFC" => data_out<= x"EA";
        when x"3DFD" => data_out<= x"EA";
        when x"3DFE" => data_out<= x"EA";
        when x"3DFF" => data_out<= x"EA";
        when x"3E00" => data_out<= x"EA";
        when x"3E01" => data_out<= x"EA";
        when x"3E02" => data_out<= x"EA";
        when x"3E03" => data_out<= x"EA";
        when x"3E04" => data_out<= x"EA";
        when x"3E05" => data_out<= x"EA";
        when x"3E06" => data_out<= x"EA";
        when x"3E07" => data_out<= x"EA";
        when x"3E08" => data_out<= x"EA";
        when x"3E09" => data_out<= x"EA";
        when x"3E0A" => data_out<= x"EA";
        when x"3E0B" => data_out<= x"EA";
        when x"3E0C" => data_out<= x"EA";
        when x"3E0D" => data_out<= x"EA";
        when x"3E0E" => data_out<= x"EA";
        when x"3E0F" => data_out<= x"EA";
        when x"3E10" => data_out<= x"EA";
        when x"3E11" => data_out<= x"EA";
        when x"3E12" => data_out<= x"EA";
        when x"3E13" => data_out<= x"EA";
        when x"3E14" => data_out<= x"EA";
        when x"3E15" => data_out<= x"EA";
        when x"3E16" => data_out<= x"EA";
        when x"3E17" => data_out<= x"EA";
        when x"3E18" => data_out<= x"EA";
        when x"3E19" => data_out<= x"EA";
        when x"3E1A" => data_out<= x"EA";
        when x"3E1B" => data_out<= x"EA";
        when x"3E1C" => data_out<= x"EA";
        when x"3E1D" => data_out<= x"EA";
        when x"3E1E" => data_out<= x"EA";
        when x"3E1F" => data_out<= x"EA";
        when x"3E20" => data_out<= x"EA";
        when x"3E21" => data_out<= x"EA";
        when x"3E22" => data_out<= x"EA";
        when x"3E23" => data_out<= x"EA";
        when x"3E24" => data_out<= x"EA";
        when x"3E25" => data_out<= x"EA";
        when x"3E26" => data_out<= x"EA";
        when x"3E27" => data_out<= x"EA";
        when x"3E28" => data_out<= x"EA";
        when x"3E29" => data_out<= x"EA";
        when x"3E2A" => data_out<= x"EA";
        when x"3E2B" => data_out<= x"EA";
        when x"3E2C" => data_out<= x"EA";
        when x"3E2D" => data_out<= x"EA";
        when x"3E2E" => data_out<= x"EA";
        when x"3E2F" => data_out<= x"EA";
        when x"3E30" => data_out<= x"EA";
        when x"3E31" => data_out<= x"EA";
        when x"3E32" => data_out<= x"EA";
        when x"3E33" => data_out<= x"EA";
        when x"3E34" => data_out<= x"EA";
        when x"3E35" => data_out<= x"EA";
        when x"3E36" => data_out<= x"EA";
        when x"3E37" => data_out<= x"EA";
        when x"3E38" => data_out<= x"EA";
        when x"3E39" => data_out<= x"EA";
        when x"3E3A" => data_out<= x"EA";
        when x"3E3B" => data_out<= x"EA";
        when x"3E3C" => data_out<= x"EA";
        when x"3E3D" => data_out<= x"EA";
        when x"3E3E" => data_out<= x"EA";
        when x"3E3F" => data_out<= x"EA";
        when x"3E40" => data_out<= x"EA";
        when x"3E41" => data_out<= x"EA";
        when x"3E42" => data_out<= x"EA";
        when x"3E43" => data_out<= x"EA";
        when x"3E44" => data_out<= x"EA";
        when x"3E45" => data_out<= x"EA";
        when x"3E46" => data_out<= x"EA";
        when x"3E47" => data_out<= x"EA";
        when x"3E48" => data_out<= x"EA";
        when x"3E49" => data_out<= x"EA";
        when x"3E4A" => data_out<= x"EA";
        when x"3E4B" => data_out<= x"EA";
        when x"3E4C" => data_out<= x"EA";
        when x"3E4D" => data_out<= x"EA";
        when x"3E4E" => data_out<= x"EA";
        when x"3E4F" => data_out<= x"EA";
        when x"3E50" => data_out<= x"EA";
        when x"3E51" => data_out<= x"EA";
        when x"3E52" => data_out<= x"EA";
        when x"3E53" => data_out<= x"EA";
        when x"3E54" => data_out<= x"EA";
        when x"3E55" => data_out<= x"EA";
        when x"3E56" => data_out<= x"EA";
        when x"3E57" => data_out<= x"EA";
        when x"3E58" => data_out<= x"EA";
        when x"3E59" => data_out<= x"EA";
        when x"3E5A" => data_out<= x"EA";
        when x"3E5B" => data_out<= x"EA";
        when x"3E5C" => data_out<= x"EA";
        when x"3E5D" => data_out<= x"EA";
        when x"3E5E" => data_out<= x"EA";
        when x"3E5F" => data_out<= x"EA";
        when x"3E60" => data_out<= x"EA";
        when x"3E61" => data_out<= x"EA";
        when x"3E62" => data_out<= x"EA";
        when x"3E63" => data_out<= x"EA";
        when x"3E64" => data_out<= x"EA";
        when x"3E65" => data_out<= x"EA";
        when x"3E66" => data_out<= x"EA";
        when x"3E67" => data_out<= x"EA";
        when x"3E68" => data_out<= x"EA";
        when x"3E69" => data_out<= x"EA";
        when x"3E6A" => data_out<= x"EA";
        when x"3E6B" => data_out<= x"EA";
        when x"3E6C" => data_out<= x"EA";
        when x"3E6D" => data_out<= x"EA";
        when x"3E6E" => data_out<= x"EA";
        when x"3E6F" => data_out<= x"EA";
        when x"3E70" => data_out<= x"EA";
        when x"3E71" => data_out<= x"EA";
        when x"3E72" => data_out<= x"EA";
        when x"3E73" => data_out<= x"EA";
        when x"3E74" => data_out<= x"EA";
        when x"3E75" => data_out<= x"EA";
        when x"3E76" => data_out<= x"EA";
        when x"3E77" => data_out<= x"EA";
        when x"3E78" => data_out<= x"EA";
        when x"3E79" => data_out<= x"EA";
        when x"3E7A" => data_out<= x"EA";
        when x"3E7B" => data_out<= x"EA";
        when x"3E7C" => data_out<= x"EA";
        when x"3E7D" => data_out<= x"EA";
        when x"3E7E" => data_out<= x"EA";
        when x"3E7F" => data_out<= x"EA";
        when x"3E80" => data_out<= x"EA";
        when x"3E81" => data_out<= x"EA";
        when x"3E82" => data_out<= x"EA";
        when x"3E83" => data_out<= x"EA";
        when x"3E84" => data_out<= x"EA";
        when x"3E85" => data_out<= x"EA";
        when x"3E86" => data_out<= x"EA";
        when x"3E87" => data_out<= x"EA";
        when x"3E88" => data_out<= x"EA";
        when x"3E89" => data_out<= x"EA";
        when x"3E8A" => data_out<= x"EA";
        when x"3E8B" => data_out<= x"EA";
        when x"3E8C" => data_out<= x"EA";
        when x"3E8D" => data_out<= x"EA";
        when x"3E8E" => data_out<= x"EA";
        when x"3E8F" => data_out<= x"EA";
        when x"3E90" => data_out<= x"EA";
        when x"3E91" => data_out<= x"EA";
        when x"3E92" => data_out<= x"EA";
        when x"3E93" => data_out<= x"EA";
        when x"3E94" => data_out<= x"EA";
        when x"3E95" => data_out<= x"EA";
        when x"3E96" => data_out<= x"EA";
        when x"3E97" => data_out<= x"EA";
        when x"3E98" => data_out<= x"EA";
        when x"3E99" => data_out<= x"EA";
        when x"3E9A" => data_out<= x"EA";
        when x"3E9B" => data_out<= x"EA";
        when x"3E9C" => data_out<= x"EA";
        when x"3E9D" => data_out<= x"EA";
        when x"3E9E" => data_out<= x"EA";
        when x"3E9F" => data_out<= x"EA";
        when x"3EA0" => data_out<= x"EA";
        when x"3EA1" => data_out<= x"EA";
        when x"3EA2" => data_out<= x"EA";
        when x"3EA3" => data_out<= x"EA";
        when x"3EA4" => data_out<= x"EA";
        when x"3EA5" => data_out<= x"EA";
        when x"3EA6" => data_out<= x"EA";
        when x"3EA7" => data_out<= x"EA";
        when x"3EA8" => data_out<= x"EA";
        when x"3EA9" => data_out<= x"EA";
        when x"3EAA" => data_out<= x"EA";
        when x"3EAB" => data_out<= x"EA";
        when x"3EAC" => data_out<= x"EA";
        when x"3EAD" => data_out<= x"EA";
        when x"3EAE" => data_out<= x"EA";
        when x"3EAF" => data_out<= x"EA";
        when x"3EB0" => data_out<= x"EA";
        when x"3EB1" => data_out<= x"EA";
        when x"3EB2" => data_out<= x"EA";
        when x"3EB3" => data_out<= x"EA";
        when x"3EB4" => data_out<= x"EA";
        when x"3EB5" => data_out<= x"EA";
        when x"3EB6" => data_out<= x"EA";
        when x"3EB7" => data_out<= x"EA";
        when x"3EB8" => data_out<= x"EA";
        when x"3EB9" => data_out<= x"EA";
        when x"3EBA" => data_out<= x"EA";
        when x"3EBB" => data_out<= x"EA";
        when x"3EBC" => data_out<= x"EA";
        when x"3EBD" => data_out<= x"EA";
        when x"3EBE" => data_out<= x"EA";
        when x"3EBF" => data_out<= x"EA";
        when x"3EC0" => data_out<= x"EA";
        when x"3EC1" => data_out<= x"EA";
        when x"3EC2" => data_out<= x"EA";
        when x"3EC3" => data_out<= x"EA";
        when x"3EC4" => data_out<= x"EA";
        when x"3EC5" => data_out<= x"EA";
        when x"3EC6" => data_out<= x"EA";
        when x"3EC7" => data_out<= x"EA";
        when x"3EC8" => data_out<= x"EA";
        when x"3EC9" => data_out<= x"EA";
        when x"3ECA" => data_out<= x"EA";
        when x"3ECB" => data_out<= x"EA";
        when x"3ECC" => data_out<= x"EA";
        when x"3ECD" => data_out<= x"EA";
        when x"3ECE" => data_out<= x"EA";
        when x"3ECF" => data_out<= x"EA";
        when x"3ED0" => data_out<= x"EA";
        when x"3ED1" => data_out<= x"EA";
        when x"3ED2" => data_out<= x"EA";
        when x"3ED3" => data_out<= x"EA";
        when x"3ED4" => data_out<= x"EA";
        when x"3ED5" => data_out<= x"EA";
        when x"3ED6" => data_out<= x"EA";
        when x"3ED7" => data_out<= x"EA";
        when x"3ED8" => data_out<= x"EA";
        when x"3ED9" => data_out<= x"EA";
        when x"3EDA" => data_out<= x"EA";
        when x"3EDB" => data_out<= x"EA";
        when x"3EDC" => data_out<= x"EA";
        when x"3EDD" => data_out<= x"EA";
        when x"3EDE" => data_out<= x"EA";
        when x"3EDF" => data_out<= x"EA";
        when x"3EE0" => data_out<= x"EA";
        when x"3EE1" => data_out<= x"EA";
        when x"3EE2" => data_out<= x"EA";
        when x"3EE3" => data_out<= x"EA";
        when x"3EE4" => data_out<= x"EA";
        when x"3EE5" => data_out<= x"EA";
        when x"3EE6" => data_out<= x"EA";
        when x"3EE7" => data_out<= x"EA";
        when x"3EE8" => data_out<= x"EA";
        when x"3EE9" => data_out<= x"EA";
        when x"3EEA" => data_out<= x"EA";
        when x"3EEB" => data_out<= x"EA";
        when x"3EEC" => data_out<= x"EA";
        when x"3EED" => data_out<= x"EA";
        when x"3EEE" => data_out<= x"EA";
        when x"3EEF" => data_out<= x"EA";
        when x"3EF0" => data_out<= x"EA";
        when x"3EF1" => data_out<= x"EA";
        when x"3EF2" => data_out<= x"EA";
        when x"3EF3" => data_out<= x"EA";
        when x"3EF4" => data_out<= x"EA";
        when x"3EF5" => data_out<= x"EA";
        when x"3EF6" => data_out<= x"EA";
        when x"3EF7" => data_out<= x"EA";
        when x"3EF8" => data_out<= x"EA";
        when x"3EF9" => data_out<= x"EA";
        when x"3EFA" => data_out<= x"EA";
        when x"3EFB" => data_out<= x"EA";
        when x"3EFC" => data_out<= x"EA";
        when x"3EFD" => data_out<= x"EA";
        when x"3EFE" => data_out<= x"EA";
        when x"3EFF" => data_out<= x"EA";
        when x"3F00" => data_out<= x"4C";
        when x"3F01" => data_out<= x"BF";
        when x"3F02" => data_out<= x"9F";
        when x"3F03" => data_out<= x"4C";
        when x"3F04" => data_out<= x"68";
        when x"3F05" => data_out<= x"A3";
        when x"3F06" => data_out<= x"4C";
        when x"3F07" => data_out<= x"E0";
        when x"3F08" => data_out<= x"A3";
        when x"3F09" => data_out<= x"4C";
        when x"3F0A" => data_out<= x"92";
        when x"3F0B" => data_out<= x"A6";
        when x"3F0C" => data_out<= x"4C";
        when x"3F0D" => data_out<= x"B9";
        when x"3F0E" => data_out<= x"A9";
        when x"3F0F" => data_out<= x"4C";
        when x"3F10" => data_out<= x"30";
        when x"3F11" => data_out<= x"AB";
        when x"3F12" => data_out<= x"4C";
        when x"3F13" => data_out<= x"51";
        when x"3F14" => data_out<= x"AA";
        when x"3F15" => data_out<= x"4C";
        when x"3F16" => data_out<= x"E5";
        when x"3F17" => data_out<= x"80";
        when x"3F18" => data_out<= x"4C";
        when x"3F19" => data_out<= x"F0";
        when x"3F1A" => data_out<= x"80";
        when x"3F1B" => data_out<= x"4C";
        when x"3F1C" => data_out<= x"FD";
        when x"3F1D" => data_out<= x"80";
        when x"3F1E" => data_out<= x"4C";
        when x"3F1F" => data_out<= x"22";
        when x"3F20" => data_out<= x"81";
        when x"3F21" => data_out<= x"4C";
        when x"3F22" => data_out<= x"0A";
        when x"3F23" => data_out<= x"81";
        when x"3F24" => data_out<= x"4C";
        when x"3F25" => data_out<= x"16";
        when x"3F26" => data_out<= x"81";
        when x"3F27" => data_out<= x"4C";
        when x"3F28" => data_out<= x"8D";
        when x"3F29" => data_out<= x"AB";
        when x"3F2A" => data_out<= x"4C";
        when x"3F2B" => data_out<= x"C7";
        when x"3F2C" => data_out<= x"AB";
        when x"3F2D" => data_out<= x"4C";
        when x"3F2E" => data_out<= x"6D";
        when x"3F2F" => data_out<= x"AD";
        when x"3F30" => data_out<= x"4C";
        when x"3F31" => data_out<= x"83";
        when x"3F32" => data_out<= x"AD";
        when x"3F33" => data_out<= x"4C";
        when x"3F34" => data_out<= x"C6";
        when x"3F35" => data_out<= x"AD";
        when x"3F36" => data_out<= x"EA";
        when x"3F37" => data_out<= x"EA";
        when x"3F38" => data_out<= x"EA";
        when x"3F39" => data_out<= x"EA";
        when x"3F3A" => data_out<= x"EA";
        when x"3F3B" => data_out<= x"EA";
        when x"3F3C" => data_out<= x"EA";
        when x"3F3D" => data_out<= x"EA";
        when x"3F3E" => data_out<= x"EA";
        when x"3F3F" => data_out<= x"EA";
        when x"3F40" => data_out<= x"EA";
        when x"3F41" => data_out<= x"EA";
        when x"3F42" => data_out<= x"EA";
        when x"3F43" => data_out<= x"EA";
        when x"3F44" => data_out<= x"EA";
        when x"3F45" => data_out<= x"EA";
        when x"3F46" => data_out<= x"EA";
        when x"3F47" => data_out<= x"EA";
        when x"3F48" => data_out<= x"EA";
        when x"3F49" => data_out<= x"EA";
        when x"3F4A" => data_out<= x"EA";
        when x"3F4B" => data_out<= x"EA";
        when x"3F4C" => data_out<= x"EA";
        when x"3F4D" => data_out<= x"EA";
        when x"3F4E" => data_out<= x"EA";
        when x"3F4F" => data_out<= x"EA";
        when x"3F50" => data_out<= x"52";
        when x"3F51" => data_out<= x"4F";
        when x"3F52" => data_out<= x"4D";
        when x"3F53" => data_out<= x"41";
        when x"3F54" => data_out<= x"50";
        when x"3F55" => data_out<= x"49";
        when x"3F56" => data_out<= x"01";
        when x"3F57" => data_out<= x"00";
        when x"3F58" => data_out<= x"EA";
        when x"3F59" => data_out<= x"EA";
        when x"3F5A" => data_out<= x"EA";
        when x"3F5B" => data_out<= x"EA";
        when x"3F5C" => data_out<= x"EA";
        when x"3F5D" => data_out<= x"EA";
        when x"3F5E" => data_out<= x"EA";
        when x"3F5F" => data_out<= x"EA";
        when x"3F60" => data_out<= x"EA";
        when x"3F61" => data_out<= x"EA";
        when x"3F62" => data_out<= x"EA";
        when x"3F63" => data_out<= x"EA";
        when x"3F64" => data_out<= x"EA";
        when x"3F65" => data_out<= x"EA";
        when x"3F66" => data_out<= x"EA";
        when x"3F67" => data_out<= x"EA";
        when x"3F68" => data_out<= x"EA";
        when x"3F69" => data_out<= x"EA";
        when x"3F6A" => data_out<= x"EA";
        when x"3F6B" => data_out<= x"EA";
        when x"3F6C" => data_out<= x"EA";
        when x"3F6D" => data_out<= x"EA";
        when x"3F6E" => data_out<= x"EA";
        when x"3F6F" => data_out<= x"EA";
        when x"3F70" => data_out<= x"EA";
        when x"3F71" => data_out<= x"EA";
        when x"3F72" => data_out<= x"EA";
        when x"3F73" => data_out<= x"EA";
        when x"3F74" => data_out<= x"EA";
        when x"3F75" => data_out<= x"EA";
        when x"3F76" => data_out<= x"EA";
        when x"3F77" => data_out<= x"EA";
        when x"3F78" => data_out<= x"EA";
        when x"3F79" => data_out<= x"EA";
        when x"3F7A" => data_out<= x"EA";
        when x"3F7B" => data_out<= x"EA";
        when x"3F7C" => data_out<= x"EA";
        when x"3F7D" => data_out<= x"EA";
        when x"3F7E" => data_out<= x"EA";
        when x"3F7F" => data_out<= x"EA";
        when x"3F80" => data_out<= x"EA";
        when x"3F81" => data_out<= x"EA";
        when x"3F82" => data_out<= x"EA";
        when x"3F83" => data_out<= x"EA";
        when x"3F84" => data_out<= x"EA";
        when x"3F85" => data_out<= x"EA";
        when x"3F86" => data_out<= x"EA";
        when x"3F87" => data_out<= x"EA";
        when x"3F88" => data_out<= x"EA";
        when x"3F89" => data_out<= x"EA";
        when x"3F8A" => data_out<= x"EA";
        when x"3F8B" => data_out<= x"EA";
        when x"3F8C" => data_out<= x"EA";
        when x"3F8D" => data_out<= x"EA";
        when x"3F8E" => data_out<= x"EA";
        when x"3F8F" => data_out<= x"EA";
        when x"3F90" => data_out<= x"EA";
        when x"3F91" => data_out<= x"EA";
        when x"3F92" => data_out<= x"EA";
        when x"3F93" => data_out<= x"EA";
        when x"3F94" => data_out<= x"EA";
        when x"3F95" => data_out<= x"EA";
        when x"3F96" => data_out<= x"EA";
        when x"3F97" => data_out<= x"EA";
        when x"3F98" => data_out<= x"EA";
        when x"3F99" => data_out<= x"EA";
        when x"3F9A" => data_out<= x"EA";
        when x"3F9B" => data_out<= x"EA";
        when x"3F9C" => data_out<= x"EA";
        when x"3F9D" => data_out<= x"EA";
        when x"3F9E" => data_out<= x"EA";
        when x"3F9F" => data_out<= x"EA";
        when x"3FA0" => data_out<= x"EA";
        when x"3FA1" => data_out<= x"EA";
        when x"3FA2" => data_out<= x"EA";
        when x"3FA3" => data_out<= x"EA";
        when x"3FA4" => data_out<= x"EA";
        when x"3FA5" => data_out<= x"EA";
        when x"3FA6" => data_out<= x"EA";
        when x"3FA7" => data_out<= x"EA";
        when x"3FA8" => data_out<= x"EA";
        when x"3FA9" => data_out<= x"EA";
        when x"3FAA" => data_out<= x"EA";
        when x"3FAB" => data_out<= x"EA";
        when x"3FAC" => data_out<= x"EA";
        when x"3FAD" => data_out<= x"EA";
        when x"3FAE" => data_out<= x"EA";
        when x"3FAF" => data_out<= x"EA";
        when x"3FB0" => data_out<= x"EA";
        when x"3FB1" => data_out<= x"EA";
        when x"3FB2" => data_out<= x"EA";
        when x"3FB3" => data_out<= x"EA";
        when x"3FB4" => data_out<= x"EA";
        when x"3FB5" => data_out<= x"EA";
        when x"3FB6" => data_out<= x"EA";
        when x"3FB7" => data_out<= x"EA";
        when x"3FB8" => data_out<= x"EA";
        when x"3FB9" => data_out<= x"EA";
        when x"3FBA" => data_out<= x"EA";
        when x"3FBB" => data_out<= x"EA";
        when x"3FBC" => data_out<= x"EA";
        when x"3FBD" => data_out<= x"EA";
        when x"3FBE" => data_out<= x"EA";
        when x"3FBF" => data_out<= x"EA";
        when x"3FC0" => data_out<= x"EA";
        when x"3FC1" => data_out<= x"EA";
        when x"3FC2" => data_out<= x"EA";
        when x"3FC3" => data_out<= x"EA";
        when x"3FC4" => data_out<= x"EA";
        when x"3FC5" => data_out<= x"EA";
        when x"3FC6" => data_out<= x"EA";
        when x"3FC7" => data_out<= x"EA";
        when x"3FC8" => data_out<= x"EA";
        when x"3FC9" => data_out<= x"EA";
        when x"3FCA" => data_out<= x"EA";
        when x"3FCB" => data_out<= x"EA";
        when x"3FCC" => data_out<= x"EA";
        when x"3FCD" => data_out<= x"EA";
        when x"3FCE" => data_out<= x"EA";
        when x"3FCF" => data_out<= x"EA";
        when x"3FD0" => data_out<= x"EA";
        when x"3FD1" => data_out<= x"EA";
        when x"3FD2" => data_out<= x"EA";
        when x"3FD3" => data_out<= x"EA";
        when x"3FD4" => data_out<= x"EA";
        when x"3FD5" => data_out<= x"EA";
        when x"3FD6" => data_out<= x"EA";
        when x"3FD7" => data_out<= x"EA";
        when x"3FD8" => data_out<= x"EA";
        when x"3FD9" => data_out<= x"EA";
        when x"3FDA" => data_out<= x"EA";
        when x"3FDB" => data_out<= x"EA";
        when x"3FDC" => data_out<= x"EA";
        when x"3FDD" => data_out<= x"EA";
        when x"3FDE" => data_out<= x"EA";
        when x"3FDF" => data_out<= x"EA";
        when x"3FE0" => data_out<= x"EA";
        when x"3FE1" => data_out<= x"EA";
        when x"3FE2" => data_out<= x"EA";
        when x"3FE3" => data_out<= x"EA";
        when x"3FE4" => data_out<= x"EA";
        when x"3FE5" => data_out<= x"EA";
        when x"3FE6" => data_out<= x"EA";
        when x"3FE7" => data_out<= x"EA";
        when x"3FE8" => data_out<= x"EA";
        when x"3FE9" => data_out<= x"EA";
        when x"3FEA" => data_out<= x"EA";
        when x"3FEB" => data_out<= x"EA";
        when x"3FEC" => data_out<= x"EA";
        when x"3FED" => data_out<= x"EA";
        when x"3FEE" => data_out<= x"EA";
        when x"3FEF" => data_out<= x"EA";
        when x"3FF0" => data_out<= x"EA";
        when x"3FF1" => data_out<= x"EA";
        when x"3FF2" => data_out<= x"EA";
        when x"3FF3" => data_out<= x"EA";
        when x"3FF4" => data_out<= x"EA";
        when x"3FF5" => data_out<= x"EA";
        when x"3FF6" => data_out<= x"EA";
        when x"3FF7" => data_out<= x"EA";
        when x"3FF8" => data_out<= x"EA";
        when x"3FF9" => data_out<= x"EA";
        when x"3FFA" => data_out<= x"E4";
        when x"3FFB" => data_out<= x"AD";
        when x"3FFC" => data_out<= x"00";
        when x"3FFD" => data_out<= x"80";
        when x"3FFE" => data_out<= x"E5";
        when x"3FFF" => data_out<= x"AD";
            when others => data_out<= x"FF";

        end case;
    end if;
	END PROCESS;
end architecture;
